-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Sun Apr 20 12:33:35 2025


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382422f",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"b7070020",
           9 => x"13060500",
          10 => x"93874707",
          11 => x"637cf600",
          12 => x"b7450000",
          13 => x"3386c740",
          14 => x"13050500",
          15 => x"938585c5",
          16 => x"ef10803e",
          17 => x"b7070020",
          18 => x"13864187",
          19 => x"9387071c",
          20 => x"637af600",
          21 => x"3386c740",
          22 => x"13854187",
          23 => x"93050000",
          24 => x"ef10c03a",
          25 => x"ef20c011",
          26 => x"b7050020",
          27 => x"93850500",
          28 => x"13060000",
          29 => x"13055000",
          30 => x"ef10004c",
          31 => x"ef10d008",
          32 => x"6f108040",
          33 => x"130101ff",
          34 => x"23261100",
          35 => x"ef10c044",
          36 => x"8320c100",
          37 => x"13051000",
          38 => x"13010101",
          39 => x"67800000",
          40 => x"130101fd",
          41 => x"b7470000",
          42 => x"232c4101",
          43 => x"130a0500",
          44 => x"1385c7a6",
          45 => x"23248102",
          46 => x"23229102",
          47 => x"23202103",
          48 => x"232e3101",
          49 => x"83244a08",
          50 => x"23261102",
          51 => x"37390000",
          52 => x"ef108042",
          53 => x"13044100",
          54 => x"93070400",
          55 => x"9309c1ff",
          56 => x"1309097f",
          57 => x"13f7f400",
          58 => x"3307e900",
          59 => x"03470700",
          60 => x"9387f7ff",
          61 => x"93d44400",
          62 => x"2384e700",
          63 => x"e39437ff",
          64 => x"13054100",
          65 => x"23060100",
          66 => x"ef10003f",
          67 => x"37450000",
          68 => x"130505a8",
          69 => x"ef10403e",
          70 => x"03278a08",
          71 => x"9377f700",
          72 => x"b307f900",
          73 => x"83c70700",
          74 => x"1304f4ff",
          75 => x"13574700",
          76 => x"2304f400",
          77 => x"e31434ff",
          78 => x"13054100",
          79 => x"ef10c03b",
          80 => x"37450000",
          81 => x"1305c5a8",
          82 => x"ef10003b",
          83 => x"8320c102",
          84 => x"03248102",
          85 => x"83244102",
          86 => x"03290102",
          87 => x"8329c101",
          88 => x"032a8101",
          89 => x"13010103",
          90 => x"67800000",
          91 => x"b70700f0",
          92 => x"03a74760",
          93 => x"93860700",
          94 => x"1377f7fe",
          95 => x"23a2e760",
          96 => x"83a74700",
          97 => x"93c71700",
          98 => x"23a2f600",
          99 => x"67800000",
         100 => x"370700f0",
         101 => x"83274700",
         102 => x"93e70720",
         103 => x"2322f700",
         104 => x"6f000000",
         105 => x"b71700f0",
         106 => x"93850700",
         107 => x"938505a0",
         108 => x"938747a0",
         109 => x"83a60700",
         110 => x"03a60500",
         111 => x"03a70700",
         112 => x"e31ad7fe",
         113 => x"b7870100",
         114 => x"b71600f0",
         115 => x"1305f0ff",
         116 => x"9387076a",
         117 => x"23a6a6a0",
         118 => x"b307f600",
         119 => x"23a4a6a0",
         120 => x"33b6c700",
         121 => x"23a4f6a0",
         122 => x"3306e600",
         123 => x"23a6c6a0",
         124 => x"370700f0",
         125 => x"83274700",
         126 => x"93c72700",
         127 => x"2322f700",
         128 => x"67800000",
         129 => x"b70700f0",
         130 => x"03a74710",
         131 => x"b70600f0",
         132 => x"93870710",
         133 => x"13778700",
         134 => x"630a0700",
         135 => x"03a74600",
         136 => x"13478700",
         137 => x"23a2e600",
         138 => x"83a78700",
         139 => x"67800000",
         140 => x"b70700f0",
         141 => x"03a74770",
         142 => x"93860700",
         143 => x"1377f7f0",
         144 => x"23a2e770",
         145 => x"83a74700",
         146 => x"93c74700",
         147 => x"23a2f600",
         148 => x"67800000",
         149 => x"b70700f0",
         150 => x"03a74740",
         151 => x"93860700",
         152 => x"137777ff",
         153 => x"23a2e740",
         154 => x"83a74700",
         155 => x"93c70701",
         156 => x"23a2f600",
         157 => x"67800000",
         158 => x"b70700f0",
         159 => x"03a74720",
         160 => x"93860700",
         161 => x"137777ff",
         162 => x"23a2e720",
         163 => x"83a74700",
         164 => x"93c70702",
         165 => x"23a2f600",
         166 => x"67800000",
         167 => x"b70700f0",
         168 => x"03a74730",
         169 => x"93860700",
         170 => x"137777ff",
         171 => x"23a2e730",
         172 => x"83a74700",
         173 => x"93c70708",
         174 => x"23a2f600",
         175 => x"67800000",
         176 => x"b70700f0",
         177 => x"23ae0700",
         178 => x"03a74700",
         179 => x"13470704",
         180 => x"23a2e700",
         181 => x"67800000",
         182 => x"b71700f0",
         183 => x"23a00790",
         184 => x"370700f0",
         185 => x"83274700",
         186 => x"93c70710",
         187 => x"2322f700",
         188 => x"67800000",
         189 => x"6f000000",
         190 => x"13050000",
         191 => x"67800000",
         192 => x"13050000",
         193 => x"67800000",
         194 => x"130101f7",
         195 => x"23221100",
         196 => x"23242100",
         197 => x"23263100",
         198 => x"23284100",
         199 => x"232a5100",
         200 => x"232c6100",
         201 => x"232e7100",
         202 => x"23208102",
         203 => x"23229102",
         204 => x"2324a102",
         205 => x"2326b102",
         206 => x"2328c102",
         207 => x"232ad102",
         208 => x"232ce102",
         209 => x"232ef102",
         210 => x"23200105",
         211 => x"23221105",
         212 => x"23242105",
         213 => x"23263105",
         214 => x"23284105",
         215 => x"232a5105",
         216 => x"232c6105",
         217 => x"232e7105",
         218 => x"23208107",
         219 => x"23229107",
         220 => x"2324a107",
         221 => x"2326b107",
         222 => x"2328c107",
         223 => x"232ad107",
         224 => x"232ce107",
         225 => x"232ef107",
         226 => x"f3222034",
         227 => x"23205108",
         228 => x"f3221034",
         229 => x"23225108",
         230 => x"83a20200",
         231 => x"23245108",
         232 => x"f3223034",
         233 => x"23265108",
         234 => x"f3272034",
         235 => x"1307b000",
         236 => x"6374f70c",
         237 => x"37070080",
         238 => x"1307d7ff",
         239 => x"b387e700",
         240 => x"13078001",
         241 => x"636ef700",
         242 => x"37470000",
         243 => x"93972700",
         244 => x"13074780",
         245 => x"b387e700",
         246 => x"83a70700",
         247 => x"67800700",
         248 => x"03258102",
         249 => x"83220108",
         250 => x"63c80200",
         251 => x"f3221034",
         252 => x"93824200",
         253 => x"73901234",
         254 => x"832fc107",
         255 => x"032f8107",
         256 => x"832e4107",
         257 => x"032e0107",
         258 => x"832dc106",
         259 => x"032d8106",
         260 => x"832c4106",
         261 => x"032c0106",
         262 => x"832bc105",
         263 => x"032b8105",
         264 => x"832a4105",
         265 => x"032a0105",
         266 => x"8329c104",
         267 => x"03298104",
         268 => x"83284104",
         269 => x"03280104",
         270 => x"8327c103",
         271 => x"03278103",
         272 => x"83264103",
         273 => x"03260103",
         274 => x"8325c102",
         275 => x"83244102",
         276 => x"03240102",
         277 => x"8323c101",
         278 => x"03238101",
         279 => x"83224101",
         280 => x"03220101",
         281 => x"8321c100",
         282 => x"03218100",
         283 => x"83204100",
         284 => x"13010109",
         285 => x"73002030",
         286 => x"93061000",
         287 => x"e3f2f6f6",
         288 => x"e360f7f6",
         289 => x"37470000",
         290 => x"93972700",
         291 => x"13078786",
         292 => x"b387e700",
         293 => x"83a70700",
         294 => x"67800700",
         295 => x"eff09fdb",
         296 => x"03258102",
         297 => x"6ff01ff4",
         298 => x"eff01fe3",
         299 => x"03258102",
         300 => x"6ff05ff3",
         301 => x"eff01fcf",
         302 => x"03258102",
         303 => x"6ff09ff2",
         304 => x"eff01fe0",
         305 => x"03258102",
         306 => x"6ff0dff1",
         307 => x"eff01fca",
         308 => x"03258102",
         309 => x"6ff01ff1",
         310 => x"eff09fd5",
         311 => x"03258102",
         312 => x"6ff05ff0",
         313 => x"eff01fd2",
         314 => x"03258102",
         315 => x"6ff09fef",
         316 => x"eff0dfda",
         317 => x"03258102",
         318 => x"6ff0dfee",
         319 => x"eff0dfd7",
         320 => x"03258102",
         321 => x"6ff01fee",
         322 => x"13050100",
         323 => x"eff05fb9",
         324 => x"03258102",
         325 => x"6ff01fed",
         326 => x"9307600d",
         327 => x"6380f81c",
         328 => x"63cc1703",
         329 => x"9307d005",
         330 => x"63c21715",
         331 => x"93078003",
         332 => x"63da1705",
         333 => x"938878fc",
         334 => x"93074002",
         335 => x"63e41705",
         336 => x"b7470000",
         337 => x"93878789",
         338 => x"93982800",
         339 => x"b388f800",
         340 => x"83a70800",
         341 => x"67800700",
         342 => x"93073019",
         343 => x"638af818",
         344 => x"938808c0",
         345 => x"9307f000",
         346 => x"63ee1701",
         347 => x"b7470000",
         348 => x"9387c792",
         349 => x"93982800",
         350 => x"b388f800",
         351 => x"83a70800",
         352 => x"67800700",
         353 => x"ef10503f",
         354 => x"93078005",
         355 => x"2320f500",
         356 => x"9307f0ff",
         357 => x"13850700",
         358 => x"6ff0dfe4",
         359 => x"b7270000",
         360 => x"23a2f500",
         361 => x"93070000",
         362 => x"13850700",
         363 => x"6ff09fe3",
         364 => x"ef10903c",
         365 => x"93079000",
         366 => x"2320f500",
         367 => x"9307f0ff",
         368 => x"13850700",
         369 => x"6ff01fe2",
         370 => x"ef10103b",
         371 => x"9307d000",
         372 => x"2320f500",
         373 => x"9307f0ff",
         374 => x"13850700",
         375 => x"6ff09fe0",
         376 => x"ef109039",
         377 => x"93072000",
         378 => x"2320f500",
         379 => x"9307f0ff",
         380 => x"13850700",
         381 => x"6ff01fdf",
         382 => x"ef101038",
         383 => x"9307f001",
         384 => x"2320f500",
         385 => x"9307f0ff",
         386 => x"13850700",
         387 => x"6ff09fdd",
         388 => x"93070000",
         389 => x"13850700",
         390 => x"6ff0dfdc",
         391 => x"13090600",
         392 => x"13840500",
         393 => x"635cc000",
         394 => x"b384c500",
         395 => x"03450400",
         396 => x"13041400",
         397 => x"eff01fa5",
         398 => x"e39a84fe",
         399 => x"13050900",
         400 => x"6ff05fda",
         401 => x"13090600",
         402 => x"13840500",
         403 => x"e358c0fe",
         404 => x"b384c500",
         405 => x"eff0dfa2",
         406 => x"2300a400",
         407 => x"13041400",
         408 => x"e39a84fe",
         409 => x"13050900",
         410 => x"6ff0dfd7",
         411 => x"9307900a",
         412 => x"e39af8f0",
         413 => x"13090000",
         414 => x"93040500",
         415 => x"13040900",
         416 => x"93090900",
         417 => x"93070900",
         418 => x"732410c8",
         419 => x"f32910c0",
         420 => x"f32710c8",
         421 => x"e31af4fe",
         422 => x"37460f00",
         423 => x"13060624",
         424 => x"93060000",
         425 => x"13850900",
         426 => x"93050400",
         427 => x"ef001018",
         428 => x"37460f00",
         429 => x"23a4a400",
         430 => x"93050400",
         431 => x"13850900",
         432 => x"13060624",
         433 => x"93060000",
         434 => x"ef008053",
         435 => x"23a0a400",
         436 => x"23a2b400",
         437 => x"13050900",
         438 => x"6ff0dfd0",
         439 => x"63120508",
         440 => x"37050020",
         441 => x"1305051c",
         442 => x"13050500",
         443 => x"6ff09fcf",
         444 => x"13090000",
         445 => x"93840500",
         446 => x"13040900",
         447 => x"93090900",
         448 => x"93070900",
         449 => x"732410c8",
         450 => x"f32910c0",
         451 => x"f32710c8",
         452 => x"e31af4fe",
         453 => x"37460f00",
         454 => x"13060624",
         455 => x"93060000",
         456 => x"13850900",
         457 => x"93050400",
         458 => x"ef005010",
         459 => x"9307803e",
         460 => x"b307f502",
         461 => x"37460f00",
         462 => x"93050400",
         463 => x"13850900",
         464 => x"13060624",
         465 => x"93060000",
         466 => x"23a4f400",
         467 => x"ef00404b",
         468 => x"23a0a400",
         469 => x"23a2b400",
         470 => x"13050900",
         471 => x"6ff09fc8",
         472 => x"b7870020",
         473 => x"93870700",
         474 => x"13070040",
         475 => x"b387e740",
         476 => x"e36cf5f6",
         477 => x"ef105020",
         478 => x"9307c000",
         479 => x"2320f500",
         480 => x"1305f0ff",
         481 => x"13050500",
         482 => x"6ff0dfc5",
         483 => x"13030500",
         484 => x"138e0500",
         485 => x"93080000",
         486 => x"63dc0500",
         487 => x"b337a000",
         488 => x"3307b040",
         489 => x"330ef740",
         490 => x"3303a040",
         491 => x"9308f0ff",
         492 => x"63dc0600",
         493 => x"b337c000",
         494 => x"b306d040",
         495 => x"93c8f8ff",
         496 => x"b386f640",
         497 => x"3306c040",
         498 => x"13070600",
         499 => x"13080300",
         500 => x"93070e00",
         501 => x"639c0628",
         502 => x"b7450000",
         503 => x"9385c596",
         504 => x"6376ce0e",
         505 => x"b7060100",
         506 => x"6378d60c",
         507 => x"93360610",
         508 => x"93b61600",
         509 => x"93963600",
         510 => x"3355d600",
         511 => x"b385a500",
         512 => x"83c50500",
         513 => x"13050002",
         514 => x"b386d500",
         515 => x"b305d540",
         516 => x"630cd500",
         517 => x"b317be00",
         518 => x"b356d300",
         519 => x"3317b600",
         520 => x"b3e7f600",
         521 => x"3318b300",
         522 => x"93550701",
         523 => x"33deb702",
         524 => x"13160701",
         525 => x"13560601",
         526 => x"b3f7b702",
         527 => x"13050e00",
         528 => x"3303c603",
         529 => x"93960701",
         530 => x"93570801",
         531 => x"b3e7d700",
         532 => x"63fe6700",
         533 => x"b307f700",
         534 => x"1305feff",
         535 => x"63e8e700",
         536 => x"63f66700",
         537 => x"1305eeff",
         538 => x"b387e700",
         539 => x"b3876740",
         540 => x"33d3b702",
         541 => x"13180801",
         542 => x"13580801",
         543 => x"b3f7b702",
         544 => x"b3066602",
         545 => x"93970701",
         546 => x"3368f800",
         547 => x"93070300",
         548 => x"637cd800",
         549 => x"33080701",
         550 => x"9307f3ff",
         551 => x"6366e800",
         552 => x"6374d800",
         553 => x"9307e3ff",
         554 => x"13150501",
         555 => x"3365f500",
         556 => x"93050000",
         557 => x"6f00000e",
         558 => x"37050001",
         559 => x"93068001",
         560 => x"e37ca6f2",
         561 => x"93060001",
         562 => x"6ff01ff3",
         563 => x"93060000",
         564 => x"630c0600",
         565 => x"b7070100",
         566 => x"637af60c",
         567 => x"93360610",
         568 => x"93b61600",
         569 => x"93963600",
         570 => x"b357d600",
         571 => x"b385f500",
         572 => x"83c70500",
         573 => x"b387d700",
         574 => x"93060002",
         575 => x"b385f640",
         576 => x"6390f60c",
         577 => x"b307ce40",
         578 => x"93051000",
         579 => x"13530701",
         580 => x"b3de6702",
         581 => x"13160701",
         582 => x"13560601",
         583 => x"93560801",
         584 => x"b3f76702",
         585 => x"13850e00",
         586 => x"330ed603",
         587 => x"93970701",
         588 => x"b3e7f600",
         589 => x"63fec701",
         590 => x"b307f700",
         591 => x"1385feff",
         592 => x"63e8e700",
         593 => x"63f6c701",
         594 => x"1385eeff",
         595 => x"b387e700",
         596 => x"b387c741",
         597 => x"33de6702",
         598 => x"13180801",
         599 => x"13580801",
         600 => x"b3f76702",
         601 => x"b306c603",
         602 => x"93970701",
         603 => x"3368f800",
         604 => x"93070e00",
         605 => x"637cd800",
         606 => x"33080701",
         607 => x"9307feff",
         608 => x"6366e800",
         609 => x"6374d800",
         610 => x"9307eeff",
         611 => x"13150501",
         612 => x"3365f500",
         613 => x"638a0800",
         614 => x"b337a000",
         615 => x"b305b040",
         616 => x"b385f540",
         617 => x"3305a040",
         618 => x"67800000",
         619 => x"b7070001",
         620 => x"93068001",
         621 => x"e37af6f2",
         622 => x"93060001",
         623 => x"6ff0dff2",
         624 => x"3317b600",
         625 => x"b356fe00",
         626 => x"13550701",
         627 => x"331ebe00",
         628 => x"b357f300",
         629 => x"b3e7c701",
         630 => x"33dea602",
         631 => x"13160701",
         632 => x"13560601",
         633 => x"3318b300",
         634 => x"b3f6a602",
         635 => x"3303c603",
         636 => x"93950601",
         637 => x"93d60701",
         638 => x"b3e6b600",
         639 => x"93050e00",
         640 => x"63fe6600",
         641 => x"b306d700",
         642 => x"9305feff",
         643 => x"63e8e600",
         644 => x"63f66600",
         645 => x"9305eeff",
         646 => x"b386e600",
         647 => x"b3866640",
         648 => x"33d3a602",
         649 => x"93970701",
         650 => x"93d70701",
         651 => x"b3f6a602",
         652 => x"33066602",
         653 => x"93960601",
         654 => x"b3e7d700",
         655 => x"93060300",
         656 => x"63fec700",
         657 => x"b307f700",
         658 => x"9306f3ff",
         659 => x"63e8e700",
         660 => x"63f6c700",
         661 => x"9306e3ff",
         662 => x"b387e700",
         663 => x"93950501",
         664 => x"b387c740",
         665 => x"b3e5d500",
         666 => x"6ff05fea",
         667 => x"6364de18",
         668 => x"b7070100",
         669 => x"63f4f604",
         670 => x"13b70610",
         671 => x"13371700",
         672 => x"13173700",
         673 => x"b7470000",
         674 => x"b3d5e600",
         675 => x"9387c796",
         676 => x"b387b700",
         677 => x"83c70700",
         678 => x"b387e700",
         679 => x"13070002",
         680 => x"b305f740",
         681 => x"6316f702",
         682 => x"13051000",
         683 => x"e3e4c6ef",
         684 => x"3335c300",
         685 => x"13351500",
         686 => x"6ff0dfed",
         687 => x"b7070001",
         688 => x"13078001",
         689 => x"e3f0f6fc",
         690 => x"13070001",
         691 => x"6ff09ffb",
         692 => x"3358f600",
         693 => x"b396b600",
         694 => x"3368d800",
         695 => x"3355fe00",
         696 => x"3317be00",
         697 => x"135e0801",
         698 => x"335fc503",
         699 => x"93160801",
         700 => x"93d60601",
         701 => x"b357f300",
         702 => x"b3e7e700",
         703 => x"13d70701",
         704 => x"3316b600",
         705 => x"3375c503",
         706 => x"b38ee603",
         707 => x"13150501",
         708 => x"3367a700",
         709 => x"13050f00",
         710 => x"637ed701",
         711 => x"3307e800",
         712 => x"1305ffff",
         713 => x"63680701",
         714 => x"6376d701",
         715 => x"1305efff",
         716 => x"33070701",
         717 => x"3307d741",
         718 => x"b35ec703",
         719 => x"93970701",
         720 => x"93d70701",
         721 => x"3377c703",
         722 => x"b386d603",
         723 => x"13170701",
         724 => x"b3e7e700",
         725 => x"13870e00",
         726 => x"63fed700",
         727 => x"b307f800",
         728 => x"1387feff",
         729 => x"63e80701",
         730 => x"63f6d700",
         731 => x"1387eeff",
         732 => x"b3870701",
         733 => x"13150501",
         734 => x"3365e500",
         735 => x"131e0601",
         736 => x"13170701",
         737 => x"13570701",
         738 => x"13580501",
         739 => x"135e0e01",
         740 => x"13560601",
         741 => x"b30ec703",
         742 => x"b387d740",
         743 => x"330ec803",
         744 => x"93d60e01",
         745 => x"3307c702",
         746 => x"3307c701",
         747 => x"3387e600",
         748 => x"3308c802",
         749 => x"6376c701",
         750 => x"b7060100",
         751 => x"3308d800",
         752 => x"93560701",
         753 => x"b3860601",
         754 => x"63e2d702",
         755 => x"e392d7ce",
         756 => x"939e0e01",
         757 => x"13170701",
         758 => x"93de0e01",
         759 => x"3313b300",
         760 => x"3307d701",
         761 => x"93050000",
         762 => x"e376e3da",
         763 => x"1305f5ff",
         764 => x"6ff01fcc",
         765 => x"93050000",
         766 => x"13050000",
         767 => x"6ff09fd9",
         768 => x"93080500",
         769 => x"13830500",
         770 => x"13070600",
         771 => x"13080500",
         772 => x"93870500",
         773 => x"63920628",
         774 => x"b7450000",
         775 => x"9385c596",
         776 => x"6376c30e",
         777 => x"b7060100",
         778 => x"6378d60c",
         779 => x"93360610",
         780 => x"93b61600",
         781 => x"93963600",
         782 => x"3355d600",
         783 => x"b385a500",
         784 => x"83c50500",
         785 => x"13050002",
         786 => x"b386d500",
         787 => x"b305d540",
         788 => x"630cd500",
         789 => x"b317b300",
         790 => x"b3d6d800",
         791 => x"3317b600",
         792 => x"b3e7f600",
         793 => x"3398b800",
         794 => x"93550701",
         795 => x"33d3b702",
         796 => x"13160701",
         797 => x"13560601",
         798 => x"b3f7b702",
         799 => x"13050300",
         800 => x"b3086602",
         801 => x"93960701",
         802 => x"93570801",
         803 => x"b3e7d700",
         804 => x"63fe1701",
         805 => x"b307f700",
         806 => x"1305f3ff",
         807 => x"63e8e700",
         808 => x"63f61701",
         809 => x"1305e3ff",
         810 => x"b387e700",
         811 => x"b3871741",
         812 => x"b3d8b702",
         813 => x"13180801",
         814 => x"13580801",
         815 => x"b3f7b702",
         816 => x"b3061603",
         817 => x"93970701",
         818 => x"3368f800",
         819 => x"93870800",
         820 => x"637cd800",
         821 => x"33080701",
         822 => x"9387f8ff",
         823 => x"6366e800",
         824 => x"6374d800",
         825 => x"9387e8ff",
         826 => x"13150501",
         827 => x"3365f500",
         828 => x"93050000",
         829 => x"67800000",
         830 => x"37050001",
         831 => x"93068001",
         832 => x"e37ca6f2",
         833 => x"93060001",
         834 => x"6ff01ff3",
         835 => x"93060000",
         836 => x"630c0600",
         837 => x"b7070100",
         838 => x"6370f60c",
         839 => x"93360610",
         840 => x"93b61600",
         841 => x"93963600",
         842 => x"b357d600",
         843 => x"b385f500",
         844 => x"83c70500",
         845 => x"b387d700",
         846 => x"93060002",
         847 => x"b385f640",
         848 => x"6396f60a",
         849 => x"b307c340",
         850 => x"93051000",
         851 => x"93580701",
         852 => x"33de1703",
         853 => x"13160701",
         854 => x"13560601",
         855 => x"93560801",
         856 => x"b3f71703",
         857 => x"13050e00",
         858 => x"3303c603",
         859 => x"93970701",
         860 => x"b3e7f600",
         861 => x"63fe6700",
         862 => x"b307f700",
         863 => x"1305feff",
         864 => x"63e8e700",
         865 => x"63f66700",
         866 => x"1305eeff",
         867 => x"b387e700",
         868 => x"b3876740",
         869 => x"33d31703",
         870 => x"13180801",
         871 => x"13580801",
         872 => x"b3f71703",
         873 => x"b3066602",
         874 => x"93970701",
         875 => x"3368f800",
         876 => x"93070300",
         877 => x"637cd800",
         878 => x"33080701",
         879 => x"9307f3ff",
         880 => x"6366e800",
         881 => x"6374d800",
         882 => x"9307e3ff",
         883 => x"13150501",
         884 => x"3365f500",
         885 => x"67800000",
         886 => x"b7070001",
         887 => x"93068001",
         888 => x"e374f6f4",
         889 => x"93060001",
         890 => x"6ff01ff4",
         891 => x"3317b600",
         892 => x"b356f300",
         893 => x"13550701",
         894 => x"3313b300",
         895 => x"b3d7f800",
         896 => x"b3e76700",
         897 => x"33d3a602",
         898 => x"13160701",
         899 => x"13560601",
         900 => x"3398b800",
         901 => x"b3f6a602",
         902 => x"b3086602",
         903 => x"93950601",
         904 => x"93d60701",
         905 => x"b3e6b600",
         906 => x"93050300",
         907 => x"63fe1601",
         908 => x"b306d700",
         909 => x"9305f3ff",
         910 => x"63e8e600",
         911 => x"63f61601",
         912 => x"9305e3ff",
         913 => x"b386e600",
         914 => x"b3861641",
         915 => x"b3d8a602",
         916 => x"93970701",
         917 => x"93d70701",
         918 => x"b3f6a602",
         919 => x"33061603",
         920 => x"93960601",
         921 => x"b3e7d700",
         922 => x"93860800",
         923 => x"63fec700",
         924 => x"b307f700",
         925 => x"9386f8ff",
         926 => x"63e8e700",
         927 => x"63f6c700",
         928 => x"9386e8ff",
         929 => x"b387e700",
         930 => x"93950501",
         931 => x"b387c740",
         932 => x"b3e5d500",
         933 => x"6ff09feb",
         934 => x"63e4d518",
         935 => x"b7070100",
         936 => x"63f4f604",
         937 => x"93b70610",
         938 => x"93b71700",
         939 => x"93973700",
         940 => x"37470000",
         941 => x"b3d5f600",
         942 => x"1307c796",
         943 => x"3307b700",
         944 => x"03470700",
         945 => x"3307f700",
         946 => x"93070002",
         947 => x"b385e740",
         948 => x"6396e702",
         949 => x"13051000",
         950 => x"e3ee66e0",
         951 => x"33b5c800",
         952 => x"13351500",
         953 => x"67800000",
         954 => x"37070001",
         955 => x"93078001",
         956 => x"e3f0e6fc",
         957 => x"93070001",
         958 => x"6ff09ffb",
         959 => x"3355e600",
         960 => x"b396b600",
         961 => x"b357e300",
         962 => x"3365d500",
         963 => x"3313b300",
         964 => x"33d7e800",
         965 => x"33676700",
         966 => x"13530501",
         967 => x"b3de6702",
         968 => x"13180501",
         969 => x"13580801",
         970 => x"93560701",
         971 => x"3316b600",
         972 => x"b3f76702",
         973 => x"330ed803",
         974 => x"93970701",
         975 => x"b3e6f600",
         976 => x"93870e00",
         977 => x"63fec601",
         978 => x"b306d500",
         979 => x"9387feff",
         980 => x"63e8a600",
         981 => x"63f6c601",
         982 => x"9387eeff",
         983 => x"b386a600",
         984 => x"b386c641",
         985 => x"33de6602",
         986 => x"13170701",
         987 => x"13570701",
         988 => x"b3f66602",
         989 => x"3308c803",
         990 => x"93960601",
         991 => x"3367d700",
         992 => x"93060e00",
         993 => x"637e0701",
         994 => x"3307e500",
         995 => x"9306feff",
         996 => x"6368a700",
         997 => x"63760701",
         998 => x"9306eeff",
         999 => x"3307a700",
        1000 => x"93970701",
        1001 => x"33e5d700",
        1002 => x"13130601",
        1003 => x"93960601",
        1004 => x"93d60601",
        1005 => x"13530301",
        1006 => x"13560601",
        1007 => x"33070741",
        1008 => x"13580501",
        1009 => x"338e6602",
        1010 => x"33036802",
        1011 => x"93570e01",
        1012 => x"b386c602",
        1013 => x"b3866600",
        1014 => x"b387d700",
        1015 => x"3308c802",
        1016 => x"63f66700",
        1017 => x"b7060100",
        1018 => x"3308d800",
        1019 => x"93d60701",
        1020 => x"b3860601",
        1021 => x"6362d702",
        1022 => x"e31cd7ce",
        1023 => x"131e0e01",
        1024 => x"93970701",
        1025 => x"135e0e01",
        1026 => x"b398b800",
        1027 => x"b387c701",
        1028 => x"93050000",
        1029 => x"e3f0f8ce",
        1030 => x"1305f5ff",
        1031 => x"6ff05fcd",
        1032 => x"93050000",
        1033 => x"13050000",
        1034 => x"67800000",
        1035 => x"13080600",
        1036 => x"93070500",
        1037 => x"13870500",
        1038 => x"63960620",
        1039 => x"b7480000",
        1040 => x"9388c896",
        1041 => x"63fcc50c",
        1042 => x"b7060100",
        1043 => x"637ed60a",
        1044 => x"93360610",
        1045 => x"93b61600",
        1046 => x"93963600",
        1047 => x"3353d600",
        1048 => x"b3886800",
        1049 => x"83c80800",
        1050 => x"13030002",
        1051 => x"b386d800",
        1052 => x"b308d340",
        1053 => x"630cd300",
        1054 => x"33971501",
        1055 => x"b356d500",
        1056 => x"33181601",
        1057 => x"33e7e600",
        1058 => x"b3171501",
        1059 => x"13560801",
        1060 => x"b356c702",
        1061 => x"13150801",
        1062 => x"13550501",
        1063 => x"3377c702",
        1064 => x"b386a602",
        1065 => x"93150701",
        1066 => x"13d70701",
        1067 => x"3367b700",
        1068 => x"637ad700",
        1069 => x"3307e800",
        1070 => x"63660701",
        1071 => x"6374d700",
        1072 => x"33070701",
        1073 => x"3307d740",
        1074 => x"b356c702",
        1075 => x"3377c702",
        1076 => x"b386a602",
        1077 => x"93970701",
        1078 => x"13170701",
        1079 => x"93d70701",
        1080 => x"b3e7e700",
        1081 => x"63fad700",
        1082 => x"b307f800",
        1083 => x"63e60701",
        1084 => x"63f4d700",
        1085 => x"b3870701",
        1086 => x"b387d740",
        1087 => x"33d51701",
        1088 => x"93050000",
        1089 => x"67800000",
        1090 => x"37030001",
        1091 => x"93068001",
        1092 => x"e37666f4",
        1093 => x"93060001",
        1094 => x"6ff05ff4",
        1095 => x"93060000",
        1096 => x"630c0600",
        1097 => x"37070100",
        1098 => x"637ee606",
        1099 => x"93360610",
        1100 => x"93b61600",
        1101 => x"93963600",
        1102 => x"3357d600",
        1103 => x"b388e800",
        1104 => x"03c70800",
        1105 => x"3307d700",
        1106 => x"93060002",
        1107 => x"b388e640",
        1108 => x"6394e606",
        1109 => x"3387c540",
        1110 => x"93550801",
        1111 => x"3356b702",
        1112 => x"13150801",
        1113 => x"13550501",
        1114 => x"93d60701",
        1115 => x"3377b702",
        1116 => x"3306a602",
        1117 => x"13170701",
        1118 => x"33e7e600",
        1119 => x"637ac700",
        1120 => x"3307e800",
        1121 => x"63660701",
        1122 => x"6374c700",
        1123 => x"33070701",
        1124 => x"3307c740",
        1125 => x"b356b702",
        1126 => x"3377b702",
        1127 => x"b386a602",
        1128 => x"6ff05ff3",
        1129 => x"37070001",
        1130 => x"93068001",
        1131 => x"e376e6f8",
        1132 => x"93060001",
        1133 => x"6ff05ff8",
        1134 => x"33181601",
        1135 => x"b3d6e500",
        1136 => x"b3171501",
        1137 => x"b3951501",
        1138 => x"3357e500",
        1139 => x"13550801",
        1140 => x"3367b700",
        1141 => x"b3d5a602",
        1142 => x"13130801",
        1143 => x"13530301",
        1144 => x"b3f6a602",
        1145 => x"b3856502",
        1146 => x"13960601",
        1147 => x"93560701",
        1148 => x"b3e6c600",
        1149 => x"63fab600",
        1150 => x"b306d800",
        1151 => x"63e60601",
        1152 => x"63f4b600",
        1153 => x"b3860601",
        1154 => x"b386b640",
        1155 => x"33d6a602",
        1156 => x"13170701",
        1157 => x"13570701",
        1158 => x"b3f6a602",
        1159 => x"33066602",
        1160 => x"93960601",
        1161 => x"3367d700",
        1162 => x"637ac700",
        1163 => x"3307e800",
        1164 => x"63660701",
        1165 => x"6374c700",
        1166 => x"33070701",
        1167 => x"3307c740",
        1168 => x"6ff09ff1",
        1169 => x"63e2d51c",
        1170 => x"37080100",
        1171 => x"63fe0605",
        1172 => x"13b80610",
        1173 => x"13381800",
        1174 => x"13183800",
        1175 => x"b7480000",
        1176 => x"33d30601",
        1177 => x"9388c896",
        1178 => x"b3886800",
        1179 => x"83c80800",
        1180 => x"13030002",
        1181 => x"b3880801",
        1182 => x"33081341",
        1183 => x"63101305",
        1184 => x"63e4b600",
        1185 => x"636cc500",
        1186 => x"3306c540",
        1187 => x"b386d540",
        1188 => x"3337c500",
        1189 => x"93070600",
        1190 => x"3387e640",
        1191 => x"13850700",
        1192 => x"93050700",
        1193 => x"67800000",
        1194 => x"b7080001",
        1195 => x"13088001",
        1196 => x"e3f616fb",
        1197 => x"13080001",
        1198 => x"6ff05ffa",
        1199 => x"b3571601",
        1200 => x"b3960601",
        1201 => x"b3e6d700",
        1202 => x"33d71501",
        1203 => x"13d30601",
        1204 => x"335f6702",
        1205 => x"139e0601",
        1206 => x"135e0e01",
        1207 => x"b3970501",
        1208 => x"b3551501",
        1209 => x"b3e5f500",
        1210 => x"93d70501",
        1211 => x"33160601",
        1212 => x"33150501",
        1213 => x"33776702",
        1214 => x"b30eee03",
        1215 => x"13170701",
        1216 => x"b3e7e700",
        1217 => x"13070f00",
        1218 => x"63fed701",
        1219 => x"b387f600",
        1220 => x"1307ffff",
        1221 => x"63e8d700",
        1222 => x"63f6d701",
        1223 => x"1307efff",
        1224 => x"b387d700",
        1225 => x"b387d741",
        1226 => x"b3de6702",
        1227 => x"93950501",
        1228 => x"93d50501",
        1229 => x"b3f76702",
        1230 => x"13830e00",
        1231 => x"330ede03",
        1232 => x"93970701",
        1233 => x"b3e5f500",
        1234 => x"63fec501",
        1235 => x"b385b600",
        1236 => x"1383feff",
        1237 => x"63e8d500",
        1238 => x"63f6c501",
        1239 => x"1383eeff",
        1240 => x"b385d500",
        1241 => x"93170701",
        1242 => x"b3e76700",
        1243 => x"b385c541",
        1244 => x"13130301",
        1245 => x"131e0601",
        1246 => x"13570601",
        1247 => x"13530301",
        1248 => x"93d70701",
        1249 => x"135e0e01",
        1250 => x"b30ec303",
        1251 => x"338ec703",
        1252 => x"3303e302",
        1253 => x"b387e702",
        1254 => x"3303c301",
        1255 => x"13d70e01",
        1256 => x"33076700",
        1257 => x"6376c701",
        1258 => x"37030100",
        1259 => x"b3876700",
        1260 => x"13530701",
        1261 => x"939e0e01",
        1262 => x"13170701",
        1263 => x"93de0e01",
        1264 => x"b307f300",
        1265 => x"3307d701",
        1266 => x"63e6f500",
        1267 => x"639ef500",
        1268 => x"637ce500",
        1269 => x"3306c740",
        1270 => x"3333c700",
        1271 => x"b306d300",
        1272 => x"13070600",
        1273 => x"b387d740",
        1274 => x"3307e540",
        1275 => x"3335e500",
        1276 => x"b385f540",
        1277 => x"b385a540",
        1278 => x"b3981501",
        1279 => x"33570701",
        1280 => x"33e5e800",
        1281 => x"b3d50501",
        1282 => x"67800000",
        1283 => x"13030500",
        1284 => x"630a0600",
        1285 => x"2300b300",
        1286 => x"1306f6ff",
        1287 => x"13031300",
        1288 => x"e31a06fe",
        1289 => x"67800000",
        1290 => x"13030500",
        1291 => x"630e0600",
        1292 => x"83830500",
        1293 => x"23007300",
        1294 => x"1306f6ff",
        1295 => x"13031300",
        1296 => x"93851500",
        1297 => x"e31606fe",
        1298 => x"67800000",
        1299 => x"630c0602",
        1300 => x"13030500",
        1301 => x"93061000",
        1302 => x"636ab500",
        1303 => x"9306f0ff",
        1304 => x"1307f6ff",
        1305 => x"3303e300",
        1306 => x"b385e500",
        1307 => x"83830500",
        1308 => x"23007300",
        1309 => x"1306f6ff",
        1310 => x"3303d300",
        1311 => x"b385d500",
        1312 => x"e31606fe",
        1313 => x"67800000",
        1314 => x"370700f0",
        1315 => x"13070710",
        1316 => x"83274700",
        1317 => x"93f78700",
        1318 => x"e38c07fe",
        1319 => x"03258700",
        1320 => x"1375f50f",
        1321 => x"67800000",
        1322 => x"f32710fc",
        1323 => x"63960700",
        1324 => x"b7f7fa02",
        1325 => x"93870708",
        1326 => x"63060500",
        1327 => x"33d5a702",
        1328 => x"1305f5ff",
        1329 => x"b70700f0",
        1330 => x"23a6a710",
        1331 => x"23a0b710",
        1332 => x"23a20710",
        1333 => x"67800000",
        1334 => x"370700f0",
        1335 => x"1375f50f",
        1336 => x"13070710",
        1337 => x"2324a700",
        1338 => x"83274700",
        1339 => x"93f70701",
        1340 => x"e38c07fe",
        1341 => x"67800000",
        1342 => x"630e0502",
        1343 => x"130101ff",
        1344 => x"23248100",
        1345 => x"23261100",
        1346 => x"13040500",
        1347 => x"03450500",
        1348 => x"630a0500",
        1349 => x"13041400",
        1350 => x"eff01ffc",
        1351 => x"03450400",
        1352 => x"e31a05fe",
        1353 => x"8320c100",
        1354 => x"03248100",
        1355 => x"13010101",
        1356 => x"67800000",
        1357 => x"67800000",
        1358 => x"130101f9",
        1359 => x"23229106",
        1360 => x"23202107",
        1361 => x"23261106",
        1362 => x"23248106",
        1363 => x"232e3105",
        1364 => x"232c4105",
        1365 => x"232a5105",
        1366 => x"23286105",
        1367 => x"23267105",
        1368 => x"23248105",
        1369 => x"23229105",
        1370 => x"13090500",
        1371 => x"93840500",
        1372 => x"f32a00fc",
        1373 => x"b7070008",
        1374 => x"232c0100",
        1375 => x"232e0100",
        1376 => x"23200102",
        1377 => x"23220102",
        1378 => x"23240102",
        1379 => x"23260102",
        1380 => x"23280102",
        1381 => x"232a0102",
        1382 => x"232c0102",
        1383 => x"232e0102",
        1384 => x"b3fafa00",
        1385 => x"732410fc",
        1386 => x"63160400",
        1387 => x"37f4fa02",
        1388 => x"13040408",
        1389 => x"97f2ffff",
        1390 => x"938242d5",
        1391 => x"73905230",
        1392 => x"37c50100",
        1393 => x"13050520",
        1394 => x"93059000",
        1395 => x"eff0dfed",
        1396 => x"b717b7d1",
        1397 => x"93879775",
        1398 => x"b337f402",
        1399 => x"93561400",
        1400 => x"37353e05",
        1401 => x"370600f0",
        1402 => x"13576400",
        1403 => x"130535d6",
        1404 => x"9386f6ff",
        1405 => x"2326d660",
        1406 => x"b725d96f",
        1407 => x"93060600",
        1408 => x"3337a702",
        1409 => x"93d7d700",
        1410 => x"13051001",
        1411 => x"2320a660",
        1412 => x"938555d8",
        1413 => x"9387f7ff",
        1414 => x"23a8f670",
        1415 => x"37260000",
        1416 => x"1306f670",
        1417 => x"23a6c670",
        1418 => x"b337b402",
        1419 => x"13576700",
        1420 => x"1307f7ff",
        1421 => x"23a0a670",
        1422 => x"93058070",
        1423 => x"13170701",
        1424 => x"23a0b640",
        1425 => x"13678700",
        1426 => x"23a0e620",
        1427 => x"1307a007",
        1428 => x"93d73701",
        1429 => x"9387f7ff",
        1430 => x"93970701",
        1431 => x"93e7c700",
        1432 => x"23a0f630",
        1433 => x"23ace600",
        1434 => x"f3224030",
        1435 => x"93e20208",
        1436 => x"73904230",
        1437 => x"f3224030",
        1438 => x"93e28200",
        1439 => x"73904230",
        1440 => x"b7220000",
        1441 => x"93828280",
        1442 => x"73900230",
        1443 => x"b7490000",
        1444 => x"1385c9a8",
        1445 => x"eff05fe6",
        1446 => x"1304f9ff",
        1447 => x"63522003",
        1448 => x"1309f0ff",
        1449 => x"03a50400",
        1450 => x"1304f4ff",
        1451 => x"93844400",
        1452 => x"eff09fe4",
        1453 => x"1385c9a8",
        1454 => x"eff01fe4",
        1455 => x"e31424ff",
        1456 => x"37450000",
        1457 => x"130505a9",
        1458 => x"eff01fe3",
        1459 => x"63960a22",
        1460 => x"b7040010",
        1461 => x"b7998888",
        1462 => x"37f4eeee",
        1463 => x"9384f4ff",
        1464 => x"93899988",
        1465 => x"1304f4ee",
        1466 => x"374a0000",
        1467 => x"b71b0000",
        1468 => x"37f9eeee",
        1469 => x"938b0b2c",
        1470 => x"1309e9ee",
        1471 => x"6f00c000",
        1472 => x"938bfbff",
        1473 => x"63860b1a",
        1474 => x"93050000",
        1475 => x"13058100",
        1476 => x"ef00d030",
        1477 => x"e31605fe",
        1478 => x"032c8100",
        1479 => x"8325c100",
        1480 => x"37160000",
        1481 => x"9357cc01",
        1482 => x"13974500",
        1483 => x"b367f700",
        1484 => x"33f79700",
        1485 => x"b3779c00",
        1486 => x"13d58501",
        1487 => x"b387e700",
        1488 => x"13d7f541",
        1489 => x"b387a700",
        1490 => x"1375d700",
        1491 => x"b387a700",
        1492 => x"33b83703",
        1493 => x"137727ff",
        1494 => x"130606e1",
        1495 => x"93060000",
        1496 => x"13050c00",
        1497 => x"938bfbff",
        1498 => x"13583800",
        1499 => x"93184800",
        1500 => x"33880841",
        1501 => x"b3870741",
        1502 => x"b387e700",
        1503 => x"13d7f741",
        1504 => x"b307fc40",
        1505 => x"3338fc00",
        1506 => x"3387e540",
        1507 => x"33070741",
        1508 => x"b3882703",
        1509 => x"33078702",
        1510 => x"33b88702",
        1511 => x"33071701",
        1512 => x"b3878702",
        1513 => x"33070701",
        1514 => x"1358f741",
        1515 => x"13783800",
        1516 => x"b307f800",
        1517 => x"33b80701",
        1518 => x"3308e800",
        1519 => x"1317e801",
        1520 => x"93d72700",
        1521 => x"b367f700",
        1522 => x"93582840",
        1523 => x"13d7c701",
        1524 => x"13934800",
        1525 => x"3367e300",
        1526 => x"33739700",
        1527 => x"33f79700",
        1528 => x"1358f841",
        1529 => x"33076700",
        1530 => x"13d38801",
        1531 => x"33076700",
        1532 => x"1373d800",
        1533 => x"33076700",
        1534 => x"33333703",
        1535 => x"137828ff",
        1536 => x"139b4700",
        1537 => x"330bfb40",
        1538 => x"131b2b00",
        1539 => x"330b6c41",
        1540 => x"13533300",
        1541 => x"131e4300",
        1542 => x"33036e40",
        1543 => x"33076740",
        1544 => x"33070701",
        1545 => x"1358f741",
        1546 => x"3387e740",
        1547 => x"33880841",
        1548 => x"b3b8e700",
        1549 => x"33081841",
        1550 => x"33032703",
        1551 => x"33088802",
        1552 => x"b3388702",
        1553 => x"33086800",
        1554 => x"33078702",
        1555 => x"33081801",
        1556 => x"9358f841",
        1557 => x"93f83800",
        1558 => x"3387e800",
        1559 => x"b3381701",
        1560 => x"b3880801",
        1561 => x"9398e801",
        1562 => x"13572700",
        1563 => x"33e7e800",
        1564 => x"13184700",
        1565 => x"3307e840",
        1566 => x"13172700",
        1567 => x"b38ce740",
        1568 => x"efe0dff0",
        1569 => x"83260101",
        1570 => x"13070500",
        1571 => x"13080b00",
        1572 => x"93870c00",
        1573 => x"13060c00",
        1574 => x"93058aaf",
        1575 => x"13058101",
        1576 => x"ef008047",
        1577 => x"13058101",
        1578 => x"eff01fc5",
        1579 => x"e39e0be4",
        1580 => x"63940a00",
        1581 => x"73001000",
        1582 => x"b70700f0",
        1583 => x"9306f00f",
        1584 => x"23a4d740",
        1585 => x"83a60720",
        1586 => x"13060009",
        1587 => x"371700f0",
        1588 => x"93e60630",
        1589 => x"23a0d720",
        1590 => x"23a4c720",
        1591 => x"83a60730",
        1592 => x"93e60630",
        1593 => x"23a0d730",
        1594 => x"23a4c730",
        1595 => x"93071000",
        1596 => x"2320f790",
        1597 => x"6ff09fdf",
        1598 => x"37450000",
        1599 => x"130505ac",
        1600 => x"eff09fbf",
        1601 => x"6ff0dfdc",
        1602 => x"130101ff",
        1603 => x"23248100",
        1604 => x"23261100",
        1605 => x"93070000",
        1606 => x"13040500",
        1607 => x"63880700",
        1608 => x"93050000",
        1609 => x"97000000",
        1610 => x"e7000000",
        1611 => x"83a74187",
        1612 => x"63840700",
        1613 => x"e7800700",
        1614 => x"13050400",
        1615 => x"ef101047",
        1616 => x"13050000",
        1617 => x"67800000",
        1618 => x"130101ff",
        1619 => x"23248100",
        1620 => x"23261100",
        1621 => x"13040500",
        1622 => x"2316b500",
        1623 => x"2317c500",
        1624 => x"23200500",
        1625 => x"23220500",
        1626 => x"23240500",
        1627 => x"23220506",
        1628 => x"23280500",
        1629 => x"232a0500",
        1630 => x"232c0500",
        1631 => x"13068000",
        1632 => x"93050000",
        1633 => x"1305c505",
        1634 => x"eff05fa8",
        1635 => x"b7270000",
        1636 => x"9387c7d8",
        1637 => x"2322f402",
        1638 => x"b7270000",
        1639 => x"938747de",
        1640 => x"2324f402",
        1641 => x"b7270000",
        1642 => x"938787e6",
        1643 => x"2326f402",
        1644 => x"b7270000",
        1645 => x"938707ec",
        1646 => x"8320c100",
        1647 => x"23208402",
        1648 => x"2328f402",
        1649 => x"03248100",
        1650 => x"13010101",
        1651 => x"67800000",
        1652 => x"b7350000",
        1653 => x"37050020",
        1654 => x"13868181",
        1655 => x"93850533",
        1656 => x"13054502",
        1657 => x"6f00c021",
        1658 => x"83254500",
        1659 => x"130101ff",
        1660 => x"b7070020",
        1661 => x"23248100",
        1662 => x"23261100",
        1663 => x"93878708",
        1664 => x"13040500",
        1665 => x"6384f500",
        1666 => x"ef109012",
        1667 => x"83258400",
        1668 => x"9387018f",
        1669 => x"6386f500",
        1670 => x"13050400",
        1671 => x"ef105011",
        1672 => x"8325c400",
        1673 => x"93878195",
        1674 => x"638cf500",
        1675 => x"13050400",
        1676 => x"03248100",
        1677 => x"8320c100",
        1678 => x"13010101",
        1679 => x"6f10500f",
        1680 => x"8320c100",
        1681 => x"03248100",
        1682 => x"13010101",
        1683 => x"67800000",
        1684 => x"b7270000",
        1685 => x"37050020",
        1686 => x"130101ff",
        1687 => x"9387079d",
        1688 => x"13060000",
        1689 => x"93054000",
        1690 => x"13058508",
        1691 => x"23261100",
        1692 => x"23aaf186",
        1693 => x"eff05fed",
        1694 => x"13061000",
        1695 => x"93059000",
        1696 => x"1385018f",
        1697 => x"eff05fec",
        1698 => x"8320c100",
        1699 => x"13062000",
        1700 => x"93052001",
        1701 => x"13858195",
        1702 => x"13010101",
        1703 => x"6ff0dfea",
        1704 => x"13050000",
        1705 => x"67800000",
        1706 => x"83a74187",
        1707 => x"130101ff",
        1708 => x"23202101",
        1709 => x"23261100",
        1710 => x"23248100",
        1711 => x"23229100",
        1712 => x"13090500",
        1713 => x"63940700",
        1714 => x"eff09ff8",
        1715 => x"93848181",
        1716 => x"03a48400",
        1717 => x"83a74400",
        1718 => x"9387f7ff",
        1719 => x"63d80702",
        1720 => x"03a40400",
        1721 => x"6310040c",
        1722 => x"9305c01a",
        1723 => x"13050900",
        1724 => x"ef00900b",
        1725 => x"13040500",
        1726 => x"63140508",
        1727 => x"23a00400",
        1728 => x"9307c000",
        1729 => x"2320f900",
        1730 => x"6f004005",
        1731 => x"0317c400",
        1732 => x"63140706",
        1733 => x"b707ffff",
        1734 => x"93871700",
        1735 => x"23220406",
        1736 => x"23200400",
        1737 => x"23220400",
        1738 => x"23240400",
        1739 => x"2326f400",
        1740 => x"23280400",
        1741 => x"232a0400",
        1742 => x"232c0400",
        1743 => x"13068000",
        1744 => x"93050000",
        1745 => x"1305c405",
        1746 => x"eff05f8c",
        1747 => x"232a0402",
        1748 => x"232c0402",
        1749 => x"23240404",
        1750 => x"23260404",
        1751 => x"8320c100",
        1752 => x"13050400",
        1753 => x"03248100",
        1754 => x"83244100",
        1755 => x"03290100",
        1756 => x"13010101",
        1757 => x"67800000",
        1758 => x"13048406",
        1759 => x"6ff0dff5",
        1760 => x"93074000",
        1761 => x"23200500",
        1762 => x"2322f500",
        1763 => x"1305c500",
        1764 => x"2324a400",
        1765 => x"1306001a",
        1766 => x"93050000",
        1767 => x"eff01f87",
        1768 => x"23a08400",
        1769 => x"93040400",
        1770 => x"6ff09ff2",
        1771 => x"83270502",
        1772 => x"639e0700",
        1773 => x"b7270000",
        1774 => x"9387879e",
        1775 => x"2320f502",
        1776 => x"83a74187",
        1777 => x"63940700",
        1778 => x"6ff09fe8",
        1779 => x"67800000",
        1780 => x"67800000",
        1781 => x"67800000",
        1782 => x"b7250000",
        1783 => x"13868181",
        1784 => x"93850594",
        1785 => x"13050000",
        1786 => x"6f008001",
        1787 => x"b7250000",
        1788 => x"13868181",
        1789 => x"938505aa",
        1790 => x"13050000",
        1791 => x"6f004000",
        1792 => x"130101fd",
        1793 => x"23248102",
        1794 => x"23202103",
        1795 => x"232e3101",
        1796 => x"232c4101",
        1797 => x"23286101",
        1798 => x"23267101",
        1799 => x"23261102",
        1800 => x"23229102",
        1801 => x"232a5101",
        1802 => x"93090500",
        1803 => x"138a0500",
        1804 => x"13040600",
        1805 => x"13090000",
        1806 => x"130b1000",
        1807 => x"930bf0ff",
        1808 => x"83248400",
        1809 => x"832a4400",
        1810 => x"938afaff",
        1811 => x"63de0a02",
        1812 => x"03240400",
        1813 => x"e31604fe",
        1814 => x"8320c102",
        1815 => x"03248102",
        1816 => x"83244102",
        1817 => x"8329c101",
        1818 => x"032a8101",
        1819 => x"832a4101",
        1820 => x"032b0101",
        1821 => x"832bc100",
        1822 => x"13050900",
        1823 => x"03290102",
        1824 => x"13010103",
        1825 => x"67800000",
        1826 => x"83d7c400",
        1827 => x"637efb00",
        1828 => x"8397e400",
        1829 => x"638a7701",
        1830 => x"93850400",
        1831 => x"13850900",
        1832 => x"e7000a00",
        1833 => x"3369a900",
        1834 => x"93848406",
        1835 => x"6ff0dff9",
        1836 => x"130101f6",
        1837 => x"232af108",
        1838 => x"b7070080",
        1839 => x"9387f7ff",
        1840 => x"232ef100",
        1841 => x"2328f100",
        1842 => x"b707ffff",
        1843 => x"2326d108",
        1844 => x"2324b100",
        1845 => x"232cb100",
        1846 => x"93878720",
        1847 => x"9306c108",
        1848 => x"93058100",
        1849 => x"232e1106",
        1850 => x"232af100",
        1851 => x"2328e108",
        1852 => x"232c0109",
        1853 => x"232e1109",
        1854 => x"23260106",
        1855 => x"2322d100",
        1856 => x"ef00103a",
        1857 => x"83278100",
        1858 => x"23800700",
        1859 => x"8320c107",
        1860 => x"1301010a",
        1861 => x"67800000",
        1862 => x"130101f6",
        1863 => x"232af108",
        1864 => x"b7070080",
        1865 => x"9387f7ff",
        1866 => x"232ef100",
        1867 => x"2328f100",
        1868 => x"b707ffff",
        1869 => x"93878720",
        1870 => x"232af100",
        1871 => x"2324a100",
        1872 => x"232ca100",
        1873 => x"03a50187",
        1874 => x"2324c108",
        1875 => x"2326d108",
        1876 => x"13860500",
        1877 => x"93068108",
        1878 => x"93058100",
        1879 => x"232e1106",
        1880 => x"2328e108",
        1881 => x"232c0109",
        1882 => x"232e1109",
        1883 => x"23260106",
        1884 => x"2322d100",
        1885 => x"ef00d032",
        1886 => x"83278100",
        1887 => x"23800700",
        1888 => x"8320c107",
        1889 => x"1301010a",
        1890 => x"67800000",
        1891 => x"130101ff",
        1892 => x"23248100",
        1893 => x"13840500",
        1894 => x"8395e500",
        1895 => x"23261100",
        1896 => x"ef008033",
        1897 => x"63400502",
        1898 => x"83274405",
        1899 => x"b387a700",
        1900 => x"232af404",
        1901 => x"8320c100",
        1902 => x"03248100",
        1903 => x"13010101",
        1904 => x"67800000",
        1905 => x"8357c400",
        1906 => x"37f7ffff",
        1907 => x"1307f7ff",
        1908 => x"b3f7e700",
        1909 => x"2316f400",
        1910 => x"6ff0dffd",
        1911 => x"13050000",
        1912 => x"67800000",
        1913 => x"83d7c500",
        1914 => x"130101fe",
        1915 => x"232c8100",
        1916 => x"232a9100",
        1917 => x"23282101",
        1918 => x"23263101",
        1919 => x"232e1100",
        1920 => x"93f70710",
        1921 => x"93040500",
        1922 => x"13840500",
        1923 => x"13090600",
        1924 => x"93890600",
        1925 => x"638a0700",
        1926 => x"8395e500",
        1927 => x"93062000",
        1928 => x"13060000",
        1929 => x"ef004026",
        1930 => x"8357c400",
        1931 => x"37f7ffff",
        1932 => x"1307f7ff",
        1933 => x"b3f7e700",
        1934 => x"8315e400",
        1935 => x"2316f400",
        1936 => x"03248101",
        1937 => x"8320c101",
        1938 => x"93860900",
        1939 => x"13060900",
        1940 => x"8329c100",
        1941 => x"03290101",
        1942 => x"13850400",
        1943 => x"83244101",
        1944 => x"13010102",
        1945 => x"6f00402c",
        1946 => x"130101ff",
        1947 => x"23248100",
        1948 => x"13840500",
        1949 => x"8395e500",
        1950 => x"23261100",
        1951 => x"ef00c020",
        1952 => x"1307f0ff",
        1953 => x"8317c400",
        1954 => x"6312e502",
        1955 => x"37f7ffff",
        1956 => x"1307f7ff",
        1957 => x"b3f7e700",
        1958 => x"2316f400",
        1959 => x"8320c100",
        1960 => x"03248100",
        1961 => x"13010101",
        1962 => x"67800000",
        1963 => x"37170000",
        1964 => x"b3e7e700",
        1965 => x"2316f400",
        1966 => x"232aa404",
        1967 => x"6ff01ffe",
        1968 => x"8395e500",
        1969 => x"6f004000",
        1970 => x"130101ff",
        1971 => x"23248100",
        1972 => x"23229100",
        1973 => x"13040500",
        1974 => x"13850500",
        1975 => x"23261100",
        1976 => x"23ac0186",
        1977 => x"ef108068",
        1978 => x"9307f0ff",
        1979 => x"6318f500",
        1980 => x"83a78187",
        1981 => x"63840700",
        1982 => x"2320f400",
        1983 => x"8320c100",
        1984 => x"03248100",
        1985 => x"83244100",
        1986 => x"13010101",
        1987 => x"67800000",
        1988 => x"83a70187",
        1989 => x"6388a716",
        1990 => x"8327c501",
        1991 => x"130101fe",
        1992 => x"232c8100",
        1993 => x"232e1100",
        1994 => x"232a9100",
        1995 => x"23282101",
        1996 => x"23263101",
        1997 => x"13040500",
        1998 => x"63840708",
        1999 => x"83a7c700",
        2000 => x"638c0702",
        2001 => x"93040000",
        2002 => x"13090008",
        2003 => x"8327c401",
        2004 => x"83a7c700",
        2005 => x"b3879700",
        2006 => x"83a50700",
        2007 => x"63980504",
        2008 => x"93844400",
        2009 => x"e39424ff",
        2010 => x"8327c401",
        2011 => x"13050400",
        2012 => x"83a5c700",
        2013 => x"ef00802b",
        2014 => x"8327c401",
        2015 => x"83a50700",
        2016 => x"63860500",
        2017 => x"13050400",
        2018 => x"ef00402a",
        2019 => x"8327c401",
        2020 => x"83a48700",
        2021 => x"63860402",
        2022 => x"93850400",
        2023 => x"13050400",
        2024 => x"83a40400",
        2025 => x"ef008028",
        2026 => x"6ff0dffe",
        2027 => x"83a90500",
        2028 => x"13050400",
        2029 => x"ef008027",
        2030 => x"93850900",
        2031 => x"6ff01ffa",
        2032 => x"83254401",
        2033 => x"63860500",
        2034 => x"13050400",
        2035 => x"ef000026",
        2036 => x"8325c401",
        2037 => x"63860500",
        2038 => x"13050400",
        2039 => x"ef000025",
        2040 => x"83250403",
        2041 => x"63860500",
        2042 => x"13050400",
        2043 => x"ef000024",
        2044 => x"83254403",
        2045 => x"63860500",
        2046 => x"13050400",
        2047 => x"ef000023",
        2048 => x"83258403",
        2049 => x"63860500",
        2050 => x"13050400",
        2051 => x"ef000022",
        2052 => x"83258404",
        2053 => x"63860500",
        2054 => x"13050400",
        2055 => x"ef000021",
        2056 => x"83254404",
        2057 => x"63860500",
        2058 => x"13050400",
        2059 => x"ef000020",
        2060 => x"8325c402",
        2061 => x"63860500",
        2062 => x"13050400",
        2063 => x"ef00001f",
        2064 => x"83270402",
        2065 => x"63820702",
        2066 => x"13050400",
        2067 => x"03248101",
        2068 => x"8320c101",
        2069 => x"83244101",
        2070 => x"03290101",
        2071 => x"8329c100",
        2072 => x"13010102",
        2073 => x"67800700",
        2074 => x"8320c101",
        2075 => x"03248101",
        2076 => x"83244101",
        2077 => x"03290101",
        2078 => x"8329c100",
        2079 => x"13010102",
        2080 => x"67800000",
        2081 => x"67800000",
        2082 => x"130101ff",
        2083 => x"23248100",
        2084 => x"23229100",
        2085 => x"13040500",
        2086 => x"13850500",
        2087 => x"93050600",
        2088 => x"13860600",
        2089 => x"23261100",
        2090 => x"23ac0186",
        2091 => x"ef10405a",
        2092 => x"9307f0ff",
        2093 => x"6318f500",
        2094 => x"83a78187",
        2095 => x"63840700",
        2096 => x"2320f400",
        2097 => x"8320c100",
        2098 => x"03248100",
        2099 => x"83244100",
        2100 => x"13010101",
        2101 => x"67800000",
        2102 => x"130101ff",
        2103 => x"23248100",
        2104 => x"23229100",
        2105 => x"13040500",
        2106 => x"13850500",
        2107 => x"93050600",
        2108 => x"13860600",
        2109 => x"23261100",
        2110 => x"23ac0186",
        2111 => x"ef104059",
        2112 => x"9307f0ff",
        2113 => x"6318f500",
        2114 => x"83a78187",
        2115 => x"63840700",
        2116 => x"2320f400",
        2117 => x"8320c100",
        2118 => x"03248100",
        2119 => x"83244100",
        2120 => x"13010101",
        2121 => x"67800000",
        2122 => x"130101ff",
        2123 => x"23248100",
        2124 => x"23229100",
        2125 => x"13040500",
        2126 => x"13850500",
        2127 => x"93050600",
        2128 => x"13860600",
        2129 => x"23261100",
        2130 => x"23ac0186",
        2131 => x"ef10c05e",
        2132 => x"9307f0ff",
        2133 => x"6318f500",
        2134 => x"83a78187",
        2135 => x"63840700",
        2136 => x"2320f400",
        2137 => x"8320c100",
        2138 => x"03248100",
        2139 => x"83244100",
        2140 => x"13010101",
        2141 => x"67800000",
        2142 => x"03a50187",
        2143 => x"67800000",
        2144 => x"130101ff",
        2145 => x"23248100",
        2146 => x"23229100",
        2147 => x"37440000",
        2148 => x"b7440000",
        2149 => x"938784c5",
        2150 => x"130484c5",
        2151 => x"3304f440",
        2152 => x"23202101",
        2153 => x"23261100",
        2154 => x"13542440",
        2155 => x"938484c5",
        2156 => x"13090000",
        2157 => x"63108904",
        2158 => x"b7440000",
        2159 => x"37440000",
        2160 => x"938784c5",
        2161 => x"130484c5",
        2162 => x"3304f440",
        2163 => x"13542440",
        2164 => x"938484c5",
        2165 => x"13090000",
        2166 => x"63188902",
        2167 => x"8320c100",
        2168 => x"03248100",
        2169 => x"83244100",
        2170 => x"03290100",
        2171 => x"13010101",
        2172 => x"67800000",
        2173 => x"83a70400",
        2174 => x"13091900",
        2175 => x"93844400",
        2176 => x"e7800700",
        2177 => x"6ff01ffb",
        2178 => x"83a70400",
        2179 => x"13091900",
        2180 => x"93844400",
        2181 => x"e7800700",
        2182 => x"6ff01ffc",
        2183 => x"13860500",
        2184 => x"93050500",
        2185 => x"03a50187",
        2186 => x"6f10c01b",
        2187 => x"638a050e",
        2188 => x"83a7c5ff",
        2189 => x"130101fe",
        2190 => x"232c8100",
        2191 => x"232e1100",
        2192 => x"1384c5ff",
        2193 => x"63d40700",
        2194 => x"3304f400",
        2195 => x"2326a100",
        2196 => x"ef004031",
        2197 => x"83a70188",
        2198 => x"0325c100",
        2199 => x"639e0700",
        2200 => x"23220400",
        2201 => x"23a08188",
        2202 => x"03248101",
        2203 => x"8320c101",
        2204 => x"13010102",
        2205 => x"6f00402f",
        2206 => x"6374f402",
        2207 => x"03260400",
        2208 => x"b306c400",
        2209 => x"639ad700",
        2210 => x"83a60700",
        2211 => x"83a74700",
        2212 => x"b386c600",
        2213 => x"2320d400",
        2214 => x"2322f400",
        2215 => x"6ff09ffc",
        2216 => x"13870700",
        2217 => x"83a74700",
        2218 => x"63840700",
        2219 => x"e37af4fe",
        2220 => x"83260700",
        2221 => x"3306d700",
        2222 => x"63188602",
        2223 => x"03260400",
        2224 => x"b386c600",
        2225 => x"2320d700",
        2226 => x"3306d700",
        2227 => x"e39ec7f8",
        2228 => x"03a60700",
        2229 => x"83a74700",
        2230 => x"b306d600",
        2231 => x"2320d700",
        2232 => x"2322f700",
        2233 => x"6ff05ff8",
        2234 => x"6378c400",
        2235 => x"9307c000",
        2236 => x"2320f500",
        2237 => x"6ff05ff7",
        2238 => x"03260400",
        2239 => x"b306c400",
        2240 => x"639ad700",
        2241 => x"83a60700",
        2242 => x"83a74700",
        2243 => x"b386c600",
        2244 => x"2320d400",
        2245 => x"2322f400",
        2246 => x"23228700",
        2247 => x"6ff0dff4",
        2248 => x"67800000",
        2249 => x"130101ff",
        2250 => x"23202101",
        2251 => x"83a7c187",
        2252 => x"23248100",
        2253 => x"23229100",
        2254 => x"23261100",
        2255 => x"93040500",
        2256 => x"13840500",
        2257 => x"63980700",
        2258 => x"93050000",
        2259 => x"ef10400e",
        2260 => x"23aea186",
        2261 => x"93050400",
        2262 => x"13850400",
        2263 => x"ef10400d",
        2264 => x"1309f0ff",
        2265 => x"63122503",
        2266 => x"1304f0ff",
        2267 => x"8320c100",
        2268 => x"13050400",
        2269 => x"03248100",
        2270 => x"83244100",
        2271 => x"03290100",
        2272 => x"13010101",
        2273 => x"67800000",
        2274 => x"13043500",
        2275 => x"1374c4ff",
        2276 => x"e30e85fc",
        2277 => x"b305a440",
        2278 => x"13850400",
        2279 => x"ef104009",
        2280 => x"e31625fd",
        2281 => x"6ff05ffc",
        2282 => x"130101fe",
        2283 => x"232a9100",
        2284 => x"93843500",
        2285 => x"93f4c4ff",
        2286 => x"23282101",
        2287 => x"232e1100",
        2288 => x"232c8100",
        2289 => x"23263101",
        2290 => x"23244101",
        2291 => x"93848400",
        2292 => x"9307c000",
        2293 => x"13090500",
        2294 => x"63fef408",
        2295 => x"93840700",
        2296 => x"63ecb408",
        2297 => x"13050900",
        2298 => x"ef00c017",
        2299 => x"83a70188",
        2300 => x"13840700",
        2301 => x"6316040a",
        2302 => x"93850400",
        2303 => x"13050900",
        2304 => x"eff05ff2",
        2305 => x"9307f0ff",
        2306 => x"13040500",
        2307 => x"6318f514",
        2308 => x"03a40188",
        2309 => x"93070400",
        2310 => x"63980710",
        2311 => x"63060412",
        2312 => x"032a0400",
        2313 => x"93050000",
        2314 => x"13050900",
        2315 => x"330a4401",
        2316 => x"ef100000",
        2317 => x"631aaa10",
        2318 => x"83270400",
        2319 => x"13050900",
        2320 => x"b384f440",
        2321 => x"93850400",
        2322 => x"eff0dfed",
        2323 => x"9307f0ff",
        2324 => x"630cf50e",
        2325 => x"83270400",
        2326 => x"b3879700",
        2327 => x"2320f400",
        2328 => x"83a70188",
        2329 => x"03a74700",
        2330 => x"6316070c",
        2331 => x"23a00188",
        2332 => x"6f000006",
        2333 => x"e3d604f6",
        2334 => x"2320f900",
        2335 => x"13050000",
        2336 => x"8320c101",
        2337 => x"03248101",
        2338 => x"83244101",
        2339 => x"03290101",
        2340 => x"8329c100",
        2341 => x"032a8100",
        2342 => x"13010102",
        2343 => x"67800000",
        2344 => x"83260400",
        2345 => x"b3869640",
        2346 => x"63ca0606",
        2347 => x"1307b000",
        2348 => x"637ad704",
        2349 => x"23209400",
        2350 => x"33079400",
        2351 => x"63908704",
        2352 => x"23a0e188",
        2353 => x"83274400",
        2354 => x"2320d700",
        2355 => x"2322f700",
        2356 => x"13050900",
        2357 => x"ef004009",
        2358 => x"1305b400",
        2359 => x"93074400",
        2360 => x"137585ff",
        2361 => x"3307f540",
        2362 => x"e30cf5f8",
        2363 => x"3304e400",
        2364 => x"b387a740",
        2365 => x"2320f400",
        2366 => x"6ff09ff8",
        2367 => x"23a2e700",
        2368 => x"6ff05ffc",
        2369 => x"03274400",
        2370 => x"63968700",
        2371 => x"23a0e188",
        2372 => x"6ff01ffc",
        2373 => x"23a2e700",
        2374 => x"6ff09ffb",
        2375 => x"93070400",
        2376 => x"03244400",
        2377 => x"6ff01fed",
        2378 => x"13840700",
        2379 => x"83a74700",
        2380 => x"6ff09fee",
        2381 => x"13870700",
        2382 => x"83a74700",
        2383 => x"e39c87fe",
        2384 => x"23220700",
        2385 => x"6ff0dff8",
        2386 => x"9307c000",
        2387 => x"2320f900",
        2388 => x"13050900",
        2389 => x"ef004001",
        2390 => x"6ff05ff2",
        2391 => x"23209500",
        2392 => x"6ff01ff7",
        2393 => x"67800000",
        2394 => x"67800000",
        2395 => x"130101fe",
        2396 => x"23282101",
        2397 => x"03a98500",
        2398 => x"232c8100",
        2399 => x"23263101",
        2400 => x"23244101",
        2401 => x"232e1100",
        2402 => x"232a9100",
        2403 => x"23225101",
        2404 => x"23206101",
        2405 => x"13840500",
        2406 => x"130a0600",
        2407 => x"93890600",
        2408 => x"63ec2613",
        2409 => x"8397c500",
        2410 => x"13070900",
        2411 => x"93f60748",
        2412 => x"638c0608",
        2413 => x"83244401",
        2414 => x"13073000",
        2415 => x"83a50501",
        2416 => x"b384e402",
        2417 => x"13072000",
        2418 => x"832a0400",
        2419 => x"130b0500",
        2420 => x"b38aba40",
        2421 => x"b3c4e402",
        2422 => x"13871900",
        2423 => x"33075701",
        2424 => x"13860400",
        2425 => x"63f6e400",
        2426 => x"93040700",
        2427 => x"13060700",
        2428 => x"93f70740",
        2429 => x"6386070a",
        2430 => x"93050600",
        2431 => x"13050b00",
        2432 => x"eff09fda",
        2433 => x"13090500",
        2434 => x"630a050a",
        2435 => x"83250401",
        2436 => x"13860a00",
        2437 => x"efe05fe1",
        2438 => x"8357c400",
        2439 => x"93f7f7b7",
        2440 => x"93e70708",
        2441 => x"2316f400",
        2442 => x"23282401",
        2443 => x"232a9400",
        2444 => x"33095901",
        2445 => x"b3845441",
        2446 => x"23202401",
        2447 => x"23249400",
        2448 => x"13890900",
        2449 => x"13870900",
        2450 => x"93090700",
        2451 => x"03250400",
        2452 => x"13860900",
        2453 => x"93050a00",
        2454 => x"efe05fdf",
        2455 => x"83278400",
        2456 => x"13050000",
        2457 => x"b3872741",
        2458 => x"2324f400",
        2459 => x"83270400",
        2460 => x"b3873701",
        2461 => x"2320f400",
        2462 => x"8320c101",
        2463 => x"03248101",
        2464 => x"83244101",
        2465 => x"03290101",
        2466 => x"8329c100",
        2467 => x"032a8100",
        2468 => x"832a4100",
        2469 => x"032b0100",
        2470 => x"13010102",
        2471 => x"67800000",
        2472 => x"13050b00",
        2473 => x"ef00505d",
        2474 => x"13090500",
        2475 => x"e31e05f6",
        2476 => x"83250401",
        2477 => x"13050b00",
        2478 => x"eff05fb7",
        2479 => x"9307c000",
        2480 => x"2320fb00",
        2481 => x"8357c400",
        2482 => x"1305f0ff",
        2483 => x"93e70704",
        2484 => x"2316f400",
        2485 => x"6ff05ffa",
        2486 => x"13890600",
        2487 => x"6ff01ff7",
        2488 => x"83278600",
        2489 => x"130101fd",
        2490 => x"232e3101",
        2491 => x"23261102",
        2492 => x"23248102",
        2493 => x"23229102",
        2494 => x"23202103",
        2495 => x"232c4101",
        2496 => x"232a5101",
        2497 => x"23286101",
        2498 => x"23267101",
        2499 => x"23248101",
        2500 => x"23229101",
        2501 => x"2320a101",
        2502 => x"93090600",
        2503 => x"63800710",
        2504 => x"832a0600",
        2505 => x"130a0500",
        2506 => x"13840500",
        2507 => x"930b3000",
        2508 => x"130c2000",
        2509 => x"03ad4a00",
        2510 => x"03ab0a00",
        2511 => x"938a8a00",
        2512 => x"e30a0dfe",
        2513 => x"03298400",
        2514 => x"93040900",
        2515 => x"63662d15",
        2516 => x"8317c400",
        2517 => x"13f70748",
        2518 => x"63060708",
        2519 => x"83244401",
        2520 => x"83250401",
        2521 => x"832c0400",
        2522 => x"b3847403",
        2523 => x"b38cbc40",
        2524 => x"13871c00",
        2525 => x"3307a701",
        2526 => x"b3c48403",
        2527 => x"13860400",
        2528 => x"63f6e400",
        2529 => x"93040700",
        2530 => x"13060700",
        2531 => x"93f70740",
        2532 => x"6386070c",
        2533 => x"93050600",
        2534 => x"13050a00",
        2535 => x"eff0dfc0",
        2536 => x"13090500",
        2537 => x"630a050c",
        2538 => x"83250401",
        2539 => x"13860c00",
        2540 => x"efe09fc7",
        2541 => x"8357c400",
        2542 => x"93f7f7b7",
        2543 => x"93e70708",
        2544 => x"2316f400",
        2545 => x"23282401",
        2546 => x"232a9400",
        2547 => x"33099901",
        2548 => x"b3849441",
        2549 => x"23202401",
        2550 => x"23249400",
        2551 => x"13090d00",
        2552 => x"93040d00",
        2553 => x"03250400",
        2554 => x"13860400",
        2555 => x"93050b00",
        2556 => x"efe0dfc5",
        2557 => x"83278400",
        2558 => x"b3872741",
        2559 => x"2324f400",
        2560 => x"83270400",
        2561 => x"b3879700",
        2562 => x"2320f400",
        2563 => x"83a78900",
        2564 => x"b387a741",
        2565 => x"23a4f900",
        2566 => x"e39e07f0",
        2567 => x"13050000",
        2568 => x"8320c102",
        2569 => x"03248102",
        2570 => x"23a20900",
        2571 => x"83244102",
        2572 => x"03290102",
        2573 => x"8329c101",
        2574 => x"032a8101",
        2575 => x"832a4101",
        2576 => x"032b0101",
        2577 => x"832bc100",
        2578 => x"032c8100",
        2579 => x"832c4100",
        2580 => x"032d0100",
        2581 => x"13010103",
        2582 => x"67800000",
        2583 => x"13050a00",
        2584 => x"ef009041",
        2585 => x"13090500",
        2586 => x"e31e05f4",
        2587 => x"83250401",
        2588 => x"13050a00",
        2589 => x"eff09f9b",
        2590 => x"9307c000",
        2591 => x"2320fa00",
        2592 => x"8357c400",
        2593 => x"1305f0ff",
        2594 => x"93e70704",
        2595 => x"2316f400",
        2596 => x"23a40900",
        2597 => x"6ff0dff8",
        2598 => x"13090d00",
        2599 => x"6ff05ff4",
        2600 => x"83d7c500",
        2601 => x"130101f6",
        2602 => x"232c8108",
        2603 => x"232a9108",
        2604 => x"23282109",
        2605 => x"23244109",
        2606 => x"232e1108",
        2607 => x"23263109",
        2608 => x"23225109",
        2609 => x"23206109",
        2610 => x"232e7107",
        2611 => x"232c8107",
        2612 => x"232a9107",
        2613 => x"93f70708",
        2614 => x"130a0500",
        2615 => x"13890500",
        2616 => x"93040600",
        2617 => x"13840600",
        2618 => x"63840706",
        2619 => x"83a70501",
        2620 => x"63900706",
        2621 => x"93050004",
        2622 => x"eff01fab",
        2623 => x"2320a900",
        2624 => x"2328a900",
        2625 => x"63120504",
        2626 => x"9307c000",
        2627 => x"2320fa00",
        2628 => x"1305f0ff",
        2629 => x"8320c109",
        2630 => x"03248109",
        2631 => x"83244109",
        2632 => x"03290109",
        2633 => x"8329c108",
        2634 => x"032a8108",
        2635 => x"832a4108",
        2636 => x"032b0108",
        2637 => x"832bc107",
        2638 => x"032c8107",
        2639 => x"832c4107",
        2640 => x"1301010a",
        2641 => x"67800000",
        2642 => x"93070004",
        2643 => x"232af900",
        2644 => x"93070002",
        2645 => x"a304f102",
        2646 => x"93070003",
        2647 => x"23220102",
        2648 => x"2305f102",
        2649 => x"23268100",
        2650 => x"930b5002",
        2651 => x"930af0ff",
        2652 => x"130c1000",
        2653 => x"130ba000",
        2654 => x"13840400",
        2655 => x"83470400",
        2656 => x"63840700",
        2657 => x"6396770d",
        2658 => x"b30c9440",
        2659 => x"63049402",
        2660 => x"93860c00",
        2661 => x"13860400",
        2662 => x"93050900",
        2663 => x"13050a00",
        2664 => x"eff0dfbc",
        2665 => x"63045525",
        2666 => x"83274102",
        2667 => x"b3879701",
        2668 => x"2322f102",
        2669 => x"83470400",
        2670 => x"638a0722",
        2671 => x"93041400",
        2672 => x"23280100",
        2673 => x"232e0100",
        2674 => x"232a5101",
        2675 => x"232c0100",
        2676 => x"a3090104",
        2677 => x"23240106",
        2678 => x"b74c0000",
        2679 => x"83c50400",
        2680 => x"13065000",
        2681 => x"13854cbc",
        2682 => x"ef00901d",
        2683 => x"03270101",
        2684 => x"93070500",
        2685 => x"13841400",
        2686 => x"63100506",
        2687 => x"93770701",
        2688 => x"63860700",
        2689 => x"93070002",
        2690 => x"a309f104",
        2691 => x"93778700",
        2692 => x"63860700",
        2693 => x"9307b002",
        2694 => x"a309f104",
        2695 => x"83c60400",
        2696 => x"9307a002",
        2697 => x"6388f604",
        2698 => x"8327c101",
        2699 => x"13840400",
        2700 => x"93060000",
        2701 => x"13069000",
        2702 => x"03470400",
        2703 => x"93051400",
        2704 => x"130707fd",
        2705 => x"637ce608",
        2706 => x"63900604",
        2707 => x"6f004005",
        2708 => x"13041400",
        2709 => x"6ff09ff2",
        2710 => x"93864cbc",
        2711 => x"b387d740",
        2712 => x"b317fc00",
        2713 => x"b3e7e700",
        2714 => x"2328f100",
        2715 => x"93040400",
        2716 => x"6ff0dff6",
        2717 => x"8327c100",
        2718 => x"93864700",
        2719 => x"83a70700",
        2720 => x"2326d100",
        2721 => x"63c60700",
        2722 => x"232ef100",
        2723 => x"6f004001",
        2724 => x"b307f040",
        2725 => x"13672700",
        2726 => x"232ef100",
        2727 => x"2328e100",
        2728 => x"03470400",
        2729 => x"9307e002",
        2730 => x"6318f706",
        2731 => x"03471400",
        2732 => x"9307a002",
        2733 => x"631ef702",
        2734 => x"8327c100",
        2735 => x"13042400",
        2736 => x"13874700",
        2737 => x"83a70700",
        2738 => x"2326e100",
        2739 => x"63d40700",
        2740 => x"9307f0ff",
        2741 => x"232af100",
        2742 => x"6f000004",
        2743 => x"b3876703",
        2744 => x"13840500",
        2745 => x"93061000",
        2746 => x"b387e700",
        2747 => x"6ff0dff4",
        2748 => x"13041400",
        2749 => x"232a0100",
        2750 => x"93060000",
        2751 => x"93070000",
        2752 => x"13069000",
        2753 => x"03470400",
        2754 => x"93051400",
        2755 => x"130707fd",
        2756 => x"6378e608",
        2757 => x"e39006fc",
        2758 => x"83450400",
        2759 => x"b7440000",
        2760 => x"13063000",
        2761 => x"1385c4bc",
        2762 => x"ef009009",
        2763 => x"63020502",
        2764 => x"83270101",
        2765 => x"9384c4bc",
        2766 => x"33059540",
        2767 => x"13070004",
        2768 => x"3317a700",
        2769 => x"b3e7e700",
        2770 => x"13041400",
        2771 => x"2328f100",
        2772 => x"83450400",
        2773 => x"37450000",
        2774 => x"13066000",
        2775 => x"130505bd",
        2776 => x"93041400",
        2777 => x"2304b102",
        2778 => x"ef009005",
        2779 => x"630a0508",
        2780 => x"93070000",
        2781 => x"63980704",
        2782 => x"03270101",
        2783 => x"8327c100",
        2784 => x"13770710",
        2785 => x"63080702",
        2786 => x"93874700",
        2787 => x"2326f100",
        2788 => x"83274102",
        2789 => x"b3873701",
        2790 => x"2322f102",
        2791 => x"6ff0dfdd",
        2792 => x"b3876703",
        2793 => x"13840500",
        2794 => x"93061000",
        2795 => x"b387e700",
        2796 => x"6ff05ff5",
        2797 => x"93877700",
        2798 => x"93f787ff",
        2799 => x"93878700",
        2800 => x"6ff0dffc",
        2801 => x"b7260000",
        2802 => x"1307c100",
        2803 => x"9386c656",
        2804 => x"13060900",
        2805 => x"93050101",
        2806 => x"13050a00",
        2807 => x"97000000",
        2808 => x"e7000000",
        2809 => x"93090500",
        2810 => x"e31455fb",
        2811 => x"8357c900",
        2812 => x"93f70704",
        2813 => x"e39e07d0",
        2814 => x"03254102",
        2815 => x"6ff09fd1",
        2816 => x"b7260000",
        2817 => x"1307c100",
        2818 => x"9386c656",
        2819 => x"13060900",
        2820 => x"93050101",
        2821 => x"13050a00",
        2822 => x"ef00c01b",
        2823 => x"6ff09ffc",
        2824 => x"130101fd",
        2825 => x"232a5101",
        2826 => x"83a70501",
        2827 => x"930a0700",
        2828 => x"03a78500",
        2829 => x"23248102",
        2830 => x"23202103",
        2831 => x"232e3101",
        2832 => x"232c4101",
        2833 => x"23261102",
        2834 => x"23229102",
        2835 => x"23286101",
        2836 => x"23267101",
        2837 => x"93090500",
        2838 => x"13840500",
        2839 => x"13090600",
        2840 => x"138a0600",
        2841 => x"63d4e700",
        2842 => x"93070700",
        2843 => x"2320f900",
        2844 => x"03473404",
        2845 => x"63060700",
        2846 => x"93871700",
        2847 => x"2320f900",
        2848 => x"83270400",
        2849 => x"93f70702",
        2850 => x"63880700",
        2851 => x"83270900",
        2852 => x"93872700",
        2853 => x"2320f900",
        2854 => x"83240400",
        2855 => x"93f46400",
        2856 => x"639e0400",
        2857 => x"130b9401",
        2858 => x"930bf0ff",
        2859 => x"8327c400",
        2860 => x"03270900",
        2861 => x"b387e740",
        2862 => x"63c4f408",
        2863 => x"83473404",
        2864 => x"b336f000",
        2865 => x"83270400",
        2866 => x"93f70702",
        2867 => x"6392070c",
        2868 => x"13063404",
        2869 => x"93050a00",
        2870 => x"13850900",
        2871 => x"e7800a00",
        2872 => x"9307f0ff",
        2873 => x"630af506",
        2874 => x"83270400",
        2875 => x"13074000",
        2876 => x"93040000",
        2877 => x"93f76700",
        2878 => x"639ee700",
        2879 => x"83270900",
        2880 => x"8324c400",
        2881 => x"b384f440",
        2882 => x"93c7f4ff",
        2883 => x"93d7f741",
        2884 => x"b3f4f400",
        2885 => x"83278400",
        2886 => x"03270401",
        2887 => x"6356f700",
        2888 => x"b387e740",
        2889 => x"b384f400",
        2890 => x"13090000",
        2891 => x"1304a401",
        2892 => x"130bf0ff",
        2893 => x"63902409",
        2894 => x"13050000",
        2895 => x"6f000002",
        2896 => x"93061000",
        2897 => x"13060b00",
        2898 => x"93050a00",
        2899 => x"13850900",
        2900 => x"e7800a00",
        2901 => x"631a7503",
        2902 => x"1305f0ff",
        2903 => x"8320c102",
        2904 => x"03248102",
        2905 => x"83244102",
        2906 => x"03290102",
        2907 => x"8329c101",
        2908 => x"032a8101",
        2909 => x"832a4101",
        2910 => x"032b0101",
        2911 => x"832bc100",
        2912 => x"13010103",
        2913 => x"67800000",
        2914 => x"93841400",
        2915 => x"6ff01ff2",
        2916 => x"3307d400",
        2917 => x"13060003",
        2918 => x"a301c704",
        2919 => x"03475404",
        2920 => x"93871600",
        2921 => x"b307f400",
        2922 => x"93862600",
        2923 => x"a381e704",
        2924 => x"6ff01ff2",
        2925 => x"93061000",
        2926 => x"13060400",
        2927 => x"93050a00",
        2928 => x"13850900",
        2929 => x"e7800a00",
        2930 => x"e30865f9",
        2931 => x"13091900",
        2932 => x"6ff05ff6",
        2933 => x"130101fd",
        2934 => x"23248102",
        2935 => x"23229102",
        2936 => x"23202103",
        2937 => x"232e3101",
        2938 => x"23261102",
        2939 => x"232c4101",
        2940 => x"232a5101",
        2941 => x"23286101",
        2942 => x"83c88501",
        2943 => x"93078007",
        2944 => x"93040500",
        2945 => x"13840500",
        2946 => x"13090600",
        2947 => x"93890600",
        2948 => x"63ee1701",
        2949 => x"93072006",
        2950 => x"93863504",
        2951 => x"63ee1701",
        2952 => x"63840828",
        2953 => x"93078005",
        2954 => x"6380f822",
        2955 => x"930a2404",
        2956 => x"23011405",
        2957 => x"6f004004",
        2958 => x"9387d8f9",
        2959 => x"93f7f70f",
        2960 => x"13065001",
        2961 => x"e364f6fe",
        2962 => x"37460000",
        2963 => x"93972700",
        2964 => x"130606c0",
        2965 => x"b387c700",
        2966 => x"83a70700",
        2967 => x"67800700",
        2968 => x"83270700",
        2969 => x"938a2504",
        2970 => x"93864700",
        2971 => x"83a70700",
        2972 => x"2320d700",
        2973 => x"2381f504",
        2974 => x"93071000",
        2975 => x"6f008026",
        2976 => x"83a70500",
        2977 => x"03250700",
        2978 => x"13f60708",
        2979 => x"93054500",
        2980 => x"63060602",
        2981 => x"83270500",
        2982 => x"2320b700",
        2983 => x"37480000",
        2984 => x"63d80700",
        2985 => x"1307d002",
        2986 => x"b307f040",
        2987 => x"a301e404",
        2988 => x"130888bd",
        2989 => x"9308a000",
        2990 => x"6f004006",
        2991 => x"13f60704",
        2992 => x"83270500",
        2993 => x"2320b700",
        2994 => x"e30a06fc",
        2995 => x"93970701",
        2996 => x"93d70741",
        2997 => x"6ff09ffc",
        2998 => x"83a50500",
        2999 => x"03260700",
        3000 => x"13f50508",
        3001 => x"83270600",
        3002 => x"13064600",
        3003 => x"631a0500",
        3004 => x"93f50504",
        3005 => x"63860500",
        3006 => x"93970701",
        3007 => x"93d70701",
        3008 => x"2320c700",
        3009 => x"37480000",
        3010 => x"1307f006",
        3011 => x"130888bd",
        3012 => x"639ae814",
        3013 => x"93088000",
        3014 => x"a3010404",
        3015 => x"03274400",
        3016 => x"2324e400",
        3017 => x"634e0700",
        3018 => x"03260400",
        3019 => x"33e7e700",
        3020 => x"938a0600",
        3021 => x"1376b6ff",
        3022 => x"2320c400",
        3023 => x"63040702",
        3024 => x"938a0600",
        3025 => x"33f71703",
        3026 => x"938afaff",
        3027 => x"3307e800",
        3028 => x"03470700",
        3029 => x"2380ea00",
        3030 => x"13870700",
        3031 => x"b3d71703",
        3032 => x"e37217ff",
        3033 => x"93078000",
        3034 => x"6394f802",
        3035 => x"83270400",
        3036 => x"93f71700",
        3037 => x"638e0700",
        3038 => x"03274400",
        3039 => x"83270401",
        3040 => x"63c8e700",
        3041 => x"93070003",
        3042 => x"a38ffafe",
        3043 => x"938afaff",
        3044 => x"b3865641",
        3045 => x"2328d400",
        3046 => x"13870900",
        3047 => x"93060900",
        3048 => x"1306c100",
        3049 => x"93050400",
        3050 => x"13850400",
        3051 => x"eff05fc7",
        3052 => x"130af0ff",
        3053 => x"631e4513",
        3054 => x"1305f0ff",
        3055 => x"8320c102",
        3056 => x"03248102",
        3057 => x"83244102",
        3058 => x"03290102",
        3059 => x"8329c101",
        3060 => x"032a8101",
        3061 => x"832a4101",
        3062 => x"032b0101",
        3063 => x"13010103",
        3064 => x"67800000",
        3065 => x"83a70500",
        3066 => x"93e70702",
        3067 => x"23a0f500",
        3068 => x"37480000",
        3069 => x"93088007",
        3070 => x"1308c8be",
        3071 => x"a3021405",
        3072 => x"03260400",
        3073 => x"83250700",
        3074 => x"13750608",
        3075 => x"83a70500",
        3076 => x"93854500",
        3077 => x"631a0500",
        3078 => x"13750604",
        3079 => x"63060500",
        3080 => x"93970701",
        3081 => x"93d70701",
        3082 => x"2320b700",
        3083 => x"13771600",
        3084 => x"63060700",
        3085 => x"13660602",
        3086 => x"2320c400",
        3087 => x"638c0700",
        3088 => x"93080001",
        3089 => x"6ff05fed",
        3090 => x"37480000",
        3091 => x"130888bd",
        3092 => x"6ff0dffa",
        3093 => x"03270400",
        3094 => x"1377f7fd",
        3095 => x"2320e400",
        3096 => x"6ff01ffe",
        3097 => x"9308a000",
        3098 => x"6ff01feb",
        3099 => x"03a60500",
        3100 => x"83270700",
        3101 => x"83a54501",
        3102 => x"13780608",
        3103 => x"13854700",
        3104 => x"630a0800",
        3105 => x"2320a700",
        3106 => x"83a70700",
        3107 => x"23a0b700",
        3108 => x"6f008001",
        3109 => x"2320a700",
        3110 => x"13760604",
        3111 => x"83a70700",
        3112 => x"e30606fe",
        3113 => x"2390b700",
        3114 => x"23280400",
        3115 => x"938a0600",
        3116 => x"6ff09fee",
        3117 => x"83270700",
        3118 => x"03a64500",
        3119 => x"93050000",
        3120 => x"93864700",
        3121 => x"2320d700",
        3122 => x"83aa0700",
        3123 => x"13850a00",
        3124 => x"ef00002f",
        3125 => x"63060500",
        3126 => x"33055541",
        3127 => x"2322a400",
        3128 => x"83274400",
        3129 => x"2328f400",
        3130 => x"a3010404",
        3131 => x"6ff0dfea",
        3132 => x"83260401",
        3133 => x"13860a00",
        3134 => x"93050900",
        3135 => x"13850400",
        3136 => x"e7800900",
        3137 => x"e30a45eb",
        3138 => x"83270400",
        3139 => x"93f72700",
        3140 => x"63940704",
        3141 => x"8327c100",
        3142 => x"0325c400",
        3143 => x"e350f5ea",
        3144 => x"13850700",
        3145 => x"6ff09fe9",
        3146 => x"93061000",
        3147 => x"13060b00",
        3148 => x"93050900",
        3149 => x"13850400",
        3150 => x"e7800900",
        3151 => x"e30e45e7",
        3152 => x"938a1a00",
        3153 => x"8327c400",
        3154 => x"0327c100",
        3155 => x"b387e740",
        3156 => x"e3ccfafc",
        3157 => x"6ff01ffc",
        3158 => x"930a0000",
        3159 => x"130b9401",
        3160 => x"6ff05ffe",
        3161 => x"8397c500",
        3162 => x"130101fe",
        3163 => x"232c8100",
        3164 => x"232a9100",
        3165 => x"232e1100",
        3166 => x"23282101",
        3167 => x"23263101",
        3168 => x"13f78700",
        3169 => x"93040500",
        3170 => x"13840500",
        3171 => x"63120712",
        3172 => x"03a74500",
        3173 => x"6346e000",
        3174 => x"03a70504",
        3175 => x"6356e010",
        3176 => x"0327c402",
        3177 => x"63020710",
        3178 => x"03a90400",
        3179 => x"93963701",
        3180 => x"23a00400",
        3181 => x"63dc060a",
        3182 => x"03264405",
        3183 => x"8357c400",
        3184 => x"93f74700",
        3185 => x"638e0700",
        3186 => x"83274400",
        3187 => x"3306f640",
        3188 => x"83274403",
        3189 => x"63860700",
        3190 => x"83270404",
        3191 => x"3306f640",
        3192 => x"8327c402",
        3193 => x"83250402",
        3194 => x"93060000",
        3195 => x"13850400",
        3196 => x"e7800700",
        3197 => x"1307f0ff",
        3198 => x"8317c400",
        3199 => x"6312e502",
        3200 => x"83a60400",
        3201 => x"1307d001",
        3202 => x"636ad70e",
        3203 => x"37074020",
        3204 => x"13071700",
        3205 => x"3357d700",
        3206 => x"13771700",
        3207 => x"6300070e",
        3208 => x"03270401",
        3209 => x"23220400",
        3210 => x"2320e400",
        3211 => x"13973701",
        3212 => x"635c0700",
        3213 => x"9307f0ff",
        3214 => x"6316f500",
        3215 => x"83a70400",
        3216 => x"63940700",
        3217 => x"232aa404",
        3218 => x"83254403",
        3219 => x"23a02401",
        3220 => x"638c0504",
        3221 => x"93074404",
        3222 => x"6386f500",
        3223 => x"13850400",
        3224 => x"efe0dffc",
        3225 => x"232a0402",
        3226 => x"6f000004",
        3227 => x"83250402",
        3228 => x"13060000",
        3229 => x"93061000",
        3230 => x"13850400",
        3231 => x"e7000700",
        3232 => x"9307f0ff",
        3233 => x"13060500",
        3234 => x"e31af5f2",
        3235 => x"83a70400",
        3236 => x"e38607f2",
        3237 => x"1307d001",
        3238 => x"6386e700",
        3239 => x"13076001",
        3240 => x"639ce704",
        3241 => x"23a02401",
        3242 => x"13050000",
        3243 => x"6f00c005",
        3244 => x"83a90501",
        3245 => x"e38a09fe",
        3246 => x"03a90500",
        3247 => x"93f73700",
        3248 => x"23a03501",
        3249 => x"33093941",
        3250 => x"13070000",
        3251 => x"63940700",
        3252 => x"03a74501",
        3253 => x"2324e400",
        3254 => x"e35820fd",
        3255 => x"83278402",
        3256 => x"83250402",
        3257 => x"93060900",
        3258 => x"13860900",
        3259 => x"13850400",
        3260 => x"e7800700",
        3261 => x"6348a002",
        3262 => x"8317c400",
        3263 => x"93e70704",
        3264 => x"2316f400",
        3265 => x"1305f0ff",
        3266 => x"8320c101",
        3267 => x"03248101",
        3268 => x"83244101",
        3269 => x"03290101",
        3270 => x"8329c100",
        3271 => x"13010102",
        3272 => x"67800000",
        3273 => x"b389a900",
        3274 => x"3309a940",
        3275 => x"6ff0dffa",
        3276 => x"83a70501",
        3277 => x"638e0704",
        3278 => x"130101fe",
        3279 => x"232c8100",
        3280 => x"232e1100",
        3281 => x"13040500",
        3282 => x"630c0500",
        3283 => x"83270502",
        3284 => x"63980700",
        3285 => x"2326b100",
        3286 => x"efe05f85",
        3287 => x"8325c100",
        3288 => x"8397c500",
        3289 => x"638c0700",
        3290 => x"13050400",
        3291 => x"03248101",
        3292 => x"8320c101",
        3293 => x"13010102",
        3294 => x"6ff0dfde",
        3295 => x"8320c101",
        3296 => x"03248101",
        3297 => x"13050000",
        3298 => x"13010102",
        3299 => x"67800000",
        3300 => x"13050000",
        3301 => x"67800000",
        3302 => x"93050500",
        3303 => x"631e0500",
        3304 => x"b7350000",
        3305 => x"37050020",
        3306 => x"13868181",
        3307 => x"93850533",
        3308 => x"13054502",
        3309 => x"6fe0df84",
        3310 => x"03a50187",
        3311 => x"6ff05ff7",
        3312 => x"93f5f50f",
        3313 => x"3306c500",
        3314 => x"6316c500",
        3315 => x"13050000",
        3316 => x"67800000",
        3317 => x"83470500",
        3318 => x"e38cb7fe",
        3319 => x"13051500",
        3320 => x"6ff09ffe",
        3321 => x"130101ff",
        3322 => x"23248100",
        3323 => x"23229100",
        3324 => x"13040500",
        3325 => x"13850500",
        3326 => x"93050600",
        3327 => x"23261100",
        3328 => x"23ac0186",
        3329 => x"ef00801d",
        3330 => x"9307f0ff",
        3331 => x"6318f500",
        3332 => x"83a78187",
        3333 => x"63840700",
        3334 => x"2320f400",
        3335 => x"8320c100",
        3336 => x"03248100",
        3337 => x"83244100",
        3338 => x"13010101",
        3339 => x"67800000",
        3340 => x"130101ff",
        3341 => x"23248100",
        3342 => x"23229100",
        3343 => x"13040500",
        3344 => x"13850500",
        3345 => x"23261100",
        3346 => x"23ac0186",
        3347 => x"ef004028",
        3348 => x"9307f0ff",
        3349 => x"6318f500",
        3350 => x"83a78187",
        3351 => x"63840700",
        3352 => x"2320f400",
        3353 => x"8320c100",
        3354 => x"03248100",
        3355 => x"83244100",
        3356 => x"13010101",
        3357 => x"67800000",
        3358 => x"130101fe",
        3359 => x"232c8100",
        3360 => x"232e1100",
        3361 => x"232a9100",
        3362 => x"23282101",
        3363 => x"23263101",
        3364 => x"23244101",
        3365 => x"13040600",
        3366 => x"63940502",
        3367 => x"03248101",
        3368 => x"8320c101",
        3369 => x"83244101",
        3370 => x"03290101",
        3371 => x"8329c100",
        3372 => x"032a8100",
        3373 => x"93050600",
        3374 => x"13010102",
        3375 => x"6fe0dfee",
        3376 => x"63180602",
        3377 => x"efe09fd6",
        3378 => x"93040000",
        3379 => x"8320c101",
        3380 => x"03248101",
        3381 => x"03290101",
        3382 => x"8329c100",
        3383 => x"032a8100",
        3384 => x"13850400",
        3385 => x"83244101",
        3386 => x"13010102",
        3387 => x"67800000",
        3388 => x"130a0500",
        3389 => x"93840500",
        3390 => x"ef008005",
        3391 => x"13090500",
        3392 => x"63668500",
        3393 => x"93571500",
        3394 => x"e3e287fc",
        3395 => x"93050400",
        3396 => x"13050a00",
        3397 => x"efe05fe9",
        3398 => x"93090500",
        3399 => x"63160500",
        3400 => x"93840900",
        3401 => x"6ff09ffa",
        3402 => x"13060400",
        3403 => x"63748900",
        3404 => x"13060900",
        3405 => x"93850400",
        3406 => x"13850900",
        3407 => x"efd0dfee",
        3408 => x"93850400",
        3409 => x"13050a00",
        3410 => x"efe05fce",
        3411 => x"6ff05ffd",
        3412 => x"83a7c5ff",
        3413 => x"1385c7ff",
        3414 => x"63d80700",
        3415 => x"b385a500",
        3416 => x"83a70500",
        3417 => x"3305f500",
        3418 => x"67800000",
        3419 => x"130101ff",
        3420 => x"23261100",
        3421 => x"23248100",
        3422 => x"93089003",
        3423 => x"73000000",
        3424 => x"13040500",
        3425 => x"635a0500",
        3426 => x"33048040",
        3427 => x"efe0dfbe",
        3428 => x"23208500",
        3429 => x"1304f0ff",
        3430 => x"8320c100",
        3431 => x"13050400",
        3432 => x"03248100",
        3433 => x"13010101",
        3434 => x"67800000",
        3435 => x"9308d005",
        3436 => x"73000000",
        3437 => x"63520502",
        3438 => x"130101ff",
        3439 => x"23248100",
        3440 => x"13040500",
        3441 => x"23261100",
        3442 => x"33048040",
        3443 => x"efe0dfba",
        3444 => x"23208500",
        3445 => x"6f000000",
        3446 => x"6f000000",
        3447 => x"130101fe",
        3448 => x"232a9100",
        3449 => x"232e1100",
        3450 => x"93040500",
        3451 => x"232c8100",
        3452 => x"93083019",
        3453 => x"13050000",
        3454 => x"93050100",
        3455 => x"73000000",
        3456 => x"13040500",
        3457 => x"635a0500",
        3458 => x"33048040",
        3459 => x"efe0dfb6",
        3460 => x"23208500",
        3461 => x"1304f0ff",
        3462 => x"83274100",
        3463 => x"03270100",
        3464 => x"8320c101",
        3465 => x"23a2f400",
        3466 => x"83278100",
        3467 => x"23a0e400",
        3468 => x"1307803e",
        3469 => x"b3c7e702",
        3470 => x"13050400",
        3471 => x"03248101",
        3472 => x"23a4f400",
        3473 => x"83244101",
        3474 => x"13010102",
        3475 => x"67800000",
        3476 => x"130101ff",
        3477 => x"23261100",
        3478 => x"23248100",
        3479 => x"9308e003",
        3480 => x"73000000",
        3481 => x"13040500",
        3482 => x"635a0500",
        3483 => x"33048040",
        3484 => x"efe09fb0",
        3485 => x"23208500",
        3486 => x"1304f0ff",
        3487 => x"8320c100",
        3488 => x"13050400",
        3489 => x"03248100",
        3490 => x"13010101",
        3491 => x"67800000",
        3492 => x"130101ff",
        3493 => x"23261100",
        3494 => x"23248100",
        3495 => x"9308f003",
        3496 => x"73000000",
        3497 => x"13040500",
        3498 => x"635a0500",
        3499 => x"33048040",
        3500 => x"efe09fac",
        3501 => x"23208500",
        3502 => x"1304f0ff",
        3503 => x"8320c100",
        3504 => x"13050400",
        3505 => x"03248100",
        3506 => x"13010101",
        3507 => x"67800000",
        3508 => x"93070500",
        3509 => x"03a54188",
        3510 => x"130101ff",
        3511 => x"23261100",
        3512 => x"631a0502",
        3513 => x"9308600d",
        3514 => x"73000000",
        3515 => x"9306f0ff",
        3516 => x"6310d502",
        3517 => x"efe05fa8",
        3518 => x"9307c000",
        3519 => x"2320f500",
        3520 => x"1305f0ff",
        3521 => x"8320c100",
        3522 => x"13010101",
        3523 => x"67800000",
        3524 => x"23a2a188",
        3525 => x"9308600d",
        3526 => x"3385a700",
        3527 => x"73000000",
        3528 => x"93060500",
        3529 => x"03a54188",
        3530 => x"b387a700",
        3531 => x"e394f6fc",
        3532 => x"23a2d188",
        3533 => x"6ff01ffd",
        3534 => x"130101ff",
        3535 => x"23261100",
        3536 => x"23248100",
        3537 => x"93080004",
        3538 => x"73000000",
        3539 => x"13040500",
        3540 => x"635a0500",
        3541 => x"33048040",
        3542 => x"efe01fa2",
        3543 => x"23208500",
        3544 => x"1304f0ff",
        3545 => x"8320c100",
        3546 => x"13050400",
        3547 => x"03248100",
        3548 => x"13010101",
        3549 => x"67800000",
        3550 => x"10000000",
        3551 => x"00000000",
        3552 => x"037a5200",
        3553 => x"017c0101",
        3554 => x"1b0c0200",
        3555 => x"10000000",
        3556 => x"18000000",
        3557 => x"f8cfffff",
        3558 => x"74040000",
        3559 => x"00000000",
        3560 => x"10000000",
        3561 => x"00000000",
        3562 => x"037a5200",
        3563 => x"017c0101",
        3564 => x"1b0c0200",
        3565 => x"10000000",
        3566 => x"18000000",
        3567 => x"44d4ffff",
        3568 => x"2c040000",
        3569 => x"00000000",
        3570 => x"10000000",
        3571 => x"00000000",
        3572 => x"037a5200",
        3573 => x"017c0101",
        3574 => x"1b0c0200",
        3575 => x"10000000",
        3576 => x"18000000",
        3577 => x"48d8ffff",
        3578 => x"e0030000",
        3579 => x"00000000",
        3580 => x"30313233",
        3581 => x"34353637",
        3582 => x"38396162",
        3583 => x"63646566",
        3584 => x"00000000",
        3585 => x"a8040000",
        3586 => x"e0030000",
        3587 => x"e0030000",
        3588 => x"e0030000",
        3589 => x"b4040000",
        3590 => x"e0030000",
        3591 => x"e0030000",
        3592 => x"e0030000",
        3593 => x"e0030000",
        3594 => x"e0030000",
        3595 => x"e0030000",
        3596 => x"e0030000",
        3597 => x"e0030000",
        3598 => x"e0030000",
        3599 => x"e0030000",
        3600 => x"c0040000",
        3601 => x"e0030000",
        3602 => x"cc040000",
        3603 => x"d8040000",
        3604 => x"e0030000",
        3605 => x"e4040000",
        3606 => x"f0040000",
        3607 => x"e0030000",
        3608 => x"fc040000",
        3609 => x"9c040000",
        3610 => x"e0030000",
        3611 => x"e0030000",
        3612 => x"e0030000",
        3613 => x"08050000",
        3614 => x"e0030000",
        3615 => x"e0030000",
        3616 => x"e0030000",
        3617 => x"e0030000",
        3618 => x"e0030000",
        3619 => x"e0030000",
        3620 => x"e0030000",
        3621 => x"18050000",
        3622 => x"b0050000",
        3623 => x"84050000",
        3624 => x"84050000",
        3625 => x"84050000",
        3626 => x"84050000",
        3627 => x"10060000",
        3628 => x"44060000",
        3629 => x"1c060000",
        3630 => x"84050000",
        3631 => x"84050000",
        3632 => x"84050000",
        3633 => x"84050000",
        3634 => x"84050000",
        3635 => x"84050000",
        3636 => x"84050000",
        3637 => x"84050000",
        3638 => x"84050000",
        3639 => x"84050000",
        3640 => x"84050000",
        3641 => x"84050000",
        3642 => x"84050000",
        3643 => x"84050000",
        3644 => x"9c050000",
        3645 => x"9c050000",
        3646 => x"84050000",
        3647 => x"84050000",
        3648 => x"84050000",
        3649 => x"84050000",
        3650 => x"84050000",
        3651 => x"84050000",
        3652 => x"84050000",
        3653 => x"84050000",
        3654 => x"84050000",
        3655 => x"84050000",
        3656 => x"84050000",
        3657 => x"84050000",
        3658 => x"10060000",
        3659 => x"b0050000",
        3660 => x"f8050000",
        3661 => x"e0050000",
        3662 => x"84050000",
        3663 => x"84050000",
        3664 => x"84050000",
        3665 => x"84050000",
        3666 => x"84050000",
        3667 => x"84050000",
        3668 => x"c8050000",
        3669 => x"84050000",
        3670 => x"84050000",
        3671 => x"84050000",
        3672 => x"84050000",
        3673 => x"9c050000",
        3674 => x"9c050000",
        3675 => x"00010202",
        3676 => x"03030303",
        3677 => x"04040404",
        3678 => x"04040404",
        3679 => x"05050505",
        3680 => x"05050505",
        3681 => x"05050505",
        3682 => x"05050505",
        3683 => x"06060606",
        3684 => x"06060606",
        3685 => x"06060606",
        3686 => x"06060606",
        3687 => x"06060606",
        3688 => x"06060606",
        3689 => x"06060606",
        3690 => x"06060606",
        3691 => x"07070707",
        3692 => x"07070707",
        3693 => x"07070707",
        3694 => x"07070707",
        3695 => x"07070707",
        3696 => x"07070707",
        3697 => x"07070707",
        3698 => x"07070707",
        3699 => x"07070707",
        3700 => x"07070707",
        3701 => x"07070707",
        3702 => x"07070707",
        3703 => x"07070707",
        3704 => x"07070707",
        3705 => x"07070707",
        3706 => x"07070707",
        3707 => x"08080808",
        3708 => x"08080808",
        3709 => x"08080808",
        3710 => x"08080808",
        3711 => x"08080808",
        3712 => x"08080808",
        3713 => x"08080808",
        3714 => x"08080808",
        3715 => x"08080808",
        3716 => x"08080808",
        3717 => x"08080808",
        3718 => x"08080808",
        3719 => x"08080808",
        3720 => x"08080808",
        3721 => x"08080808",
        3722 => x"08080808",
        3723 => x"08080808",
        3724 => x"08080808",
        3725 => x"08080808",
        3726 => x"08080808",
        3727 => x"08080808",
        3728 => x"08080808",
        3729 => x"08080808",
        3730 => x"08080808",
        3731 => x"08080808",
        3732 => x"08080808",
        3733 => x"08080808",
        3734 => x"08080808",
        3735 => x"08080808",
        3736 => x"08080808",
        3737 => x"08080808",
        3738 => x"08080808",
        3739 => x"0d0a4542",
        3740 => x"5245414b",
        3741 => x"21206d65",
        3742 => x"7063203d",
        3743 => x"20000000",
        3744 => x"20696e73",
        3745 => x"6e203d20",
        3746 => x"00000000",
        3747 => x"0d0a0000",
        3748 => x"0d0a0a44",
        3749 => x"6973706c",
        3750 => x"6179696e",
        3751 => x"67207468",
        3752 => x"65207469",
        3753 => x"6d652070",
        3754 => x"61737365",
        3755 => x"64207369",
        3756 => x"6e636520",
        3757 => x"72657365",
        3758 => x"740d0a0a",
        3759 => x"00000000",
        3760 => x"4f6e2d63",
        3761 => x"68697020",
        3762 => x"64656275",
        3763 => x"67676572",
        3764 => x"20666f75",
        3765 => x"6e642c20",
        3766 => x"736b6970",
        3767 => x"70696e67",
        3768 => x"20454252",
        3769 => x"45414b20",
        3770 => x"696e7374",
        3771 => x"72756374",
        3772 => x"696f6e0d",
        3773 => x"0a0d0a00",
        3774 => x"2530356c",
        3775 => x"643a2530",
        3776 => x"366c6420",
        3777 => x"20202530",
        3778 => x"326c643a",
        3779 => x"2530326c",
        3780 => x"643a2530",
        3781 => x"326c640d",
        3782 => x"00000000",
        3783 => x"696e7465",
        3784 => x"72727570",
        3785 => x"745f6469",
        3786 => x"72656374",
        3787 => x"00000000",
        3788 => x"54485541",
        3789 => x"53205249",
        3790 => x"53432d56",
        3791 => x"20525633",
        3792 => x"32494d20",
        3793 => x"62617265",
        3794 => x"206d6574",
        3795 => x"616c2070",
        3796 => x"726f6365",
        3797 => x"73736f72",
        3798 => x"00000000",
        3799 => x"54686520",
        3800 => x"48616775",
        3801 => x"6520556e",
        3802 => x"69766572",
        3803 => x"73697479",
        3804 => x"206f6620",
        3805 => x"4170706c",
        3806 => x"69656420",
        3807 => x"53636965",
        3808 => x"6e636573",
        3809 => x"00000000",
        3810 => x"44657061",
        3811 => x"72746d65",
        3812 => x"6e74206f",
        3813 => x"6620456c",
        3814 => x"65637472",
        3815 => x"6963616c",
        3816 => x"20456e67",
        3817 => x"696e6565",
        3818 => x"72696e67",
        3819 => x"00000000",
        3820 => x"4a2e452e",
        3821 => x"4a2e206f",
        3822 => x"70206465",
        3823 => x"6e204272",
        3824 => x"6f757700",
        3825 => x"232d302b",
        3826 => x"20000000",
        3827 => x"686c4c00",
        3828 => x"65666745",
        3829 => x"46470000",
        3830 => x"30313233",
        3831 => x"34353637",
        3832 => x"38394142",
        3833 => x"43444546",
        3834 => x"00000000",
        3835 => x"30313233",
        3836 => x"34353637",
        3837 => x"38396162",
        3838 => x"63646566",
        3839 => x"00000000",
        3840 => x"602e0000",
        3841 => x"802e0000",
        3842 => x"2c2e0000",
        3843 => x"2c2e0000",
        3844 => x"2c2e0000",
        3845 => x"2c2e0000",
        3846 => x"802e0000",
        3847 => x"2c2e0000",
        3848 => x"2c2e0000",
        3849 => x"2c2e0000",
        3850 => x"2c2e0000",
        3851 => x"6c300000",
        3852 => x"d82e0000",
        3853 => x"e42f0000",
        3854 => x"2c2e0000",
        3855 => x"2c2e0000",
        3856 => x"b4300000",
        3857 => x"2c2e0000",
        3858 => x"d82e0000",
        3859 => x"2c2e0000",
        3860 => x"2c2e0000",
        3861 => x"f02f0000",
        3862 => x"1c3b0000",
        3863 => x"303b0000",
        3864 => x"5c3b0000",
        3865 => x"883b0000",
        3866 => x"b03b0000",
        3867 => x"00000000",
        3868 => x"00000000",
        3869 => x"03000000",
        3870 => x"88000020",
        3871 => x"00000000",
        3872 => x"88000020",
        3873 => x"f0000020",
        3874 => x"58010020",
        3875 => x"00000000",
        3876 => x"00000000",
        3877 => x"00000000",
        3878 => x"00000000",
        3879 => x"00000000",
        3880 => x"00000000",
        3881 => x"00000000",
        3882 => x"00000000",
        3883 => x"00000000",
        3884 => x"00000000",
        3885 => x"00000000",
        3886 => x"00000000",
        3887 => x"00000000",
        3888 => x"00000000",
        3889 => x"00000000",
        3890 => x"24000020"
            );
end package rom_image;
