-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Sun Nov 23 17:20:28 2025


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382022f",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"37060020",
           9 => x"13050500",
          10 => x"13064607",
          11 => x"637ac500",
          12 => x"b7450000",
          13 => x"3306a640",
          14 => x"938545d8",
          15 => x"ef100039",
          16 => x"37060020",
          17 => x"13854187",
          18 => x"1306061c",
          19 => x"6378c500",
          20 => x"3306a640",
          21 => x"93050000",
          22 => x"ef108035",
          23 => x"ef20c027",
          24 => x"b7050020",
          25 => x"93850500",
          26 => x"13060000",
          27 => x"13055000",
          28 => x"ef10405f",
          29 => x"ef10501f",
          30 => x"6f10403b",
          31 => x"130101fe",
          32 => x"232e1100",
          33 => x"2326a100",
          34 => x"ef10403f",
          35 => x"8320c101",
          36 => x"0325c100",
          37 => x"13010102",
          38 => x"67800000",
          39 => x"130101fd",
          40 => x"b7470000",
          41 => x"232c4101",
          42 => x"130a0500",
          43 => x"1385c7b6",
          44 => x"23248102",
          45 => x"23229102",
          46 => x"23202103",
          47 => x"232e3101",
          48 => x"83244a08",
          49 => x"23261102",
          50 => x"37490000",
          51 => x"ef10003d",
          52 => x"13044100",
          53 => x"93070400",
          54 => x"9309c1ff",
          55 => x"13090992",
          56 => x"13f7f400",
          57 => x"3307e900",
          58 => x"03470700",
          59 => x"9387f7ff",
          60 => x"93d44400",
          61 => x"2384e700",
          62 => x"e39437ff",
          63 => x"13054100",
          64 => x"23060100",
          65 => x"ef108039",
          66 => x"37450000",
          67 => x"130505b8",
          68 => x"ef10c038",
          69 => x"03278a08",
          70 => x"9377f700",
          71 => x"b307f900",
          72 => x"83c70700",
          73 => x"1304f4ff",
          74 => x"13574700",
          75 => x"2304f400",
          76 => x"e31434ff",
          77 => x"13054100",
          78 => x"ef104036",
          79 => x"37450000",
          80 => x"1305c5b8",
          81 => x"ef108035",
          82 => x"8320c102",
          83 => x"03248102",
          84 => x"83244102",
          85 => x"03290102",
          86 => x"8329c101",
          87 => x"032a8101",
          88 => x"13010103",
          89 => x"67800000",
          90 => x"b70700f0",
          91 => x"03a74760",
          92 => x"93860700",
          93 => x"1377f7fe",
          94 => x"23a2e760",
          95 => x"83a74700",
          96 => x"93c71700",
          97 => x"23a2f600",
          98 => x"67800000",
          99 => x"370700f0",
         100 => x"83274700",
         101 => x"93e70720",
         102 => x"2322f700",
         103 => x"6f000000",
         104 => x"b71700f0",
         105 => x"b71500f0",
         106 => x"938747a0",
         107 => x"938505a0",
         108 => x"83a60700",
         109 => x"03a60500",
         110 => x"03a70700",
         111 => x"e31ad7fe",
         112 => x"b7870100",
         113 => x"b71600f0",
         114 => x"1305f0ff",
         115 => x"9387076a",
         116 => x"23a6a6a0",
         117 => x"b307f600",
         118 => x"23a4a6a0",
         119 => x"33b6c700",
         120 => x"23a4f6a0",
         121 => x"3306e600",
         122 => x"23a6c6a0",
         123 => x"370700f0",
         124 => x"83274700",
         125 => x"93c72700",
         126 => x"2322f700",
         127 => x"67800000",
         128 => x"b70700f0",
         129 => x"03a74710",
         130 => x"b70600f0",
         131 => x"93870710",
         132 => x"13778700",
         133 => x"630a0700",
         134 => x"03a74600",
         135 => x"13478700",
         136 => x"23a2e600",
         137 => x"83a78700",
         138 => x"67800000",
         139 => x"b70700f0",
         140 => x"03a74770",
         141 => x"93860700",
         142 => x"1377f7f0",
         143 => x"23a2e770",
         144 => x"83a74700",
         145 => x"93c74700",
         146 => x"23a2f600",
         147 => x"67800000",
         148 => x"b70700f0",
         149 => x"03a74740",
         150 => x"93860700",
         151 => x"137777ff",
         152 => x"23a2e740",
         153 => x"83a74700",
         154 => x"93c70701",
         155 => x"23a2f600",
         156 => x"67800000",
         157 => x"b70700f0",
         158 => x"03a74720",
         159 => x"93860700",
         160 => x"137777ff",
         161 => x"23a2e720",
         162 => x"83a74700",
         163 => x"93c70702",
         164 => x"23a2f600",
         165 => x"67800000",
         166 => x"b70700f0",
         167 => x"03a74730",
         168 => x"93860700",
         169 => x"137777ff",
         170 => x"23a2e730",
         171 => x"83a74700",
         172 => x"93c70708",
         173 => x"23a2f600",
         174 => x"67800000",
         175 => x"b70700f0",
         176 => x"23ae0700",
         177 => x"03a74700",
         178 => x"13470704",
         179 => x"23a2e700",
         180 => x"67800000",
         181 => x"b71700f0",
         182 => x"23a00790",
         183 => x"370700f0",
         184 => x"83274700",
         185 => x"93c70710",
         186 => x"2322f700",
         187 => x"67800000",
         188 => x"6f000000",
         189 => x"13050000",
         190 => x"67800000",
         191 => x"13050000",
         192 => x"67800000",
         193 => x"130101f7",
         194 => x"23221100",
         195 => x"23242100",
         196 => x"23263100",
         197 => x"23284100",
         198 => x"232a5100",
         199 => x"232c6100",
         200 => x"232e7100",
         201 => x"23208102",
         202 => x"23229102",
         203 => x"2324a102",
         204 => x"2326b102",
         205 => x"2328c102",
         206 => x"232ad102",
         207 => x"232ce102",
         208 => x"232ef102",
         209 => x"23200105",
         210 => x"23221105",
         211 => x"23242105",
         212 => x"23263105",
         213 => x"23284105",
         214 => x"232a5105",
         215 => x"232c6105",
         216 => x"232e7105",
         217 => x"23208107",
         218 => x"23229107",
         219 => x"2324a107",
         220 => x"2326b107",
         221 => x"2328c107",
         222 => x"232ad107",
         223 => x"232ce107",
         224 => x"232ef107",
         225 => x"f3222034",
         226 => x"23205108",
         227 => x"f3221034",
         228 => x"23225108",
         229 => x"83a20200",
         230 => x"23245108",
         231 => x"f3223034",
         232 => x"23265108",
         233 => x"13080100",
         234 => x"ef00400a",
         235 => x"83220108",
         236 => x"63c80200",
         237 => x"73231034",
         238 => x"13034300",
         239 => x"73101334",
         240 => x"1303b000",
         241 => x"63846200",
         242 => x"03258102",
         243 => x"832fc107",
         244 => x"032f8107",
         245 => x"832e4107",
         246 => x"032e0107",
         247 => x"832dc106",
         248 => x"032d8106",
         249 => x"832c4106",
         250 => x"032c0106",
         251 => x"832bc105",
         252 => x"032b8105",
         253 => x"832a4105",
         254 => x"032a0105",
         255 => x"8329c104",
         256 => x"03298104",
         257 => x"83284104",
         258 => x"03280104",
         259 => x"8327c103",
         260 => x"03278103",
         261 => x"83264103",
         262 => x"03260103",
         263 => x"8325c102",
         264 => x"83244102",
         265 => x"03240102",
         266 => x"8323c101",
         267 => x"03238101",
         268 => x"83224101",
         269 => x"03220101",
         270 => x"8321c100",
         271 => x"03218100",
         272 => x"83204100",
         273 => x"13010109",
         274 => x"73002030",
         275 => x"f3272034",
         276 => x"37070080",
         277 => x"1307b701",
         278 => x"6360f720",
         279 => x"130101fe",
         280 => x"37070080",
         281 => x"232e1100",
         282 => x"13072700",
         283 => x"138e0500",
         284 => x"6374f704",
         285 => x"37070080",
         286 => x"1307d7ff",
         287 => x"b387e700",
         288 => x"13078001",
         289 => x"6360f702",
         290 => x"37470000",
         291 => x"93972700",
         292 => x"13074793",
         293 => x"b387e700",
         294 => x"83a70700",
         295 => x"67800700",
         296 => x"eff05fe3",
         297 => x"13060000",
         298 => x"8320c101",
         299 => x"13050600",
         300 => x"13010102",
         301 => x"67800000",
         302 => x"13073000",
         303 => x"6386e704",
         304 => x"1307b000",
         305 => x"e390e7fe",
         306 => x"9307600d",
         307 => x"638af820",
         308 => x"63e21709",
         309 => x"9307d005",
         310 => x"63e61719",
         311 => x"93078003",
         312 => x"63f0170b",
         313 => x"938878fc",
         314 => x"93074002",
         315 => x"63ea1709",
         316 => x"b7470000",
         317 => x"93878799",
         318 => x"93982800",
         319 => x"b388f800",
         320 => x"83a70800",
         321 => x"67800700",
         322 => x"13050800",
         323 => x"eff01fb9",
         324 => x"6ff05ff9",
         325 => x"eff0dfc8",
         326 => x"6ff0dff8",
         327 => x"eff01fda",
         328 => x"6ff05ff8",
         329 => x"eff01fd5",
         330 => x"6ff0dff7",
         331 => x"eff05fd2",
         332 => x"6ff05ff7",
         333 => x"eff05fc3",
         334 => x"6ff0dff6",
         335 => x"eff01fcf",
         336 => x"6ff05ff6",
         337 => x"eff0dfcb",
         338 => x"6ff0dff5",
         339 => x"eff0dfd4",
         340 => x"6ff05ff5",
         341 => x"93073019",
         342 => x"638cf818",
         343 => x"938808c0",
         344 => x"9307f000",
         345 => x"63ee1701",
         346 => x"b7470000",
         347 => x"9387c7a2",
         348 => x"93982800",
         349 => x"b388f800",
         350 => x"83a70800",
         351 => x"67800700",
         352 => x"ef101055",
         353 => x"93078005",
         354 => x"2320f500",
         355 => x"1306f0ff",
         356 => x"6ff09ff1",
         357 => x"b7270000",
         358 => x"2322fe00",
         359 => x"6ff09ff0",
         360 => x"ef101053",
         361 => x"93079000",
         362 => x"2320f500",
         363 => x"1306f0ff",
         364 => x"6ff09fef",
         365 => x"ef10d051",
         366 => x"9307f001",
         367 => x"2320f500",
         368 => x"1306f0ff",
         369 => x"6ff05fee",
         370 => x"ef109050",
         371 => x"9307d000",
         372 => x"2320f500",
         373 => x"1306f0ff",
         374 => x"6ff01fed",
         375 => x"ef10504f",
         376 => x"93072000",
         377 => x"2320f500",
         378 => x"1306f0ff",
         379 => x"6ff0dfeb",
         380 => x"e35cc0ea",
         381 => x"232c8100",
         382 => x"3384c500",
         383 => x"03450e00",
         384 => x"130e1e00",
         385 => x"2324c100",
         386 => x"2322c101",
         387 => x"eff01fa7",
         388 => x"032e4100",
         389 => x"03268100",
         390 => x"e3128efe",
         391 => x"03248101",
         392 => x"6ff09fe8",
         393 => x"e352c0e8",
         394 => x"232c8100",
         395 => x"3384c500",
         396 => x"2324c100",
         397 => x"2322c101",
         398 => x"eff01fa4",
         399 => x"032e4100",
         400 => x"03268100",
         401 => x"2300ae00",
         402 => x"130e1e00",
         403 => x"e3128efe",
         404 => x"03248101",
         405 => x"6ff05fe5",
         406 => x"13060000",
         407 => x"13050600",
         408 => x"67800000",
         409 => x"9307900a",
         410 => x"e39cf8f0",
         411 => x"93070000",
         412 => x"2326a100",
         413 => x"13870700",
         414 => x"93860700",
         415 => x"f32710c8",
         416 => x"732710c0",
         417 => x"f32610c8",
         418 => x"e39ad7fe",
         419 => x"37460f00",
         420 => x"13060624",
         421 => x"93060000",
         422 => x"13050700",
         423 => x"93850700",
         424 => x"2324e100",
         425 => x"2322f100",
         426 => x"ef00d00e",
         427 => x"0323c100",
         428 => x"83254100",
         429 => x"37460f00",
         430 => x"2324a300",
         431 => x"03258100",
         432 => x"13060624",
         433 => x"93060000",
         434 => x"23226100",
         435 => x"ef00c04d",
         436 => x"03234100",
         437 => x"2320a300",
         438 => x"2322b300",
         439 => x"6ff09fdc",
         440 => x"63160508",
         441 => x"37060020",
         442 => x"1306061c",
         443 => x"6ff0dfdb",
         444 => x"93070000",
         445 => x"2326b100",
         446 => x"13880700",
         447 => x"13870700",
         448 => x"f32710c8",
         449 => x"732810c0",
         450 => x"732710c8",
         451 => x"e39ae7fe",
         452 => x"37460f00",
         453 => x"13060624",
         454 => x"93060000",
         455 => x"13050800",
         456 => x"93850700",
         457 => x"23240101",
         458 => x"2322f100",
         459 => x"ef009006",
         460 => x"1307803e",
         461 => x"3307e502",
         462 => x"032ec100",
         463 => x"83254100",
         464 => x"03258100",
         465 => x"37460f00",
         466 => x"13060624",
         467 => x"93060000",
         468 => x"2322c101",
         469 => x"2324ee00",
         470 => x"ef000045",
         471 => x"032e4100",
         472 => x"2320ae00",
         473 => x"2322be00",
         474 => x"6ff0dfd3",
         475 => x"b7870020",
         476 => x"93870700",
         477 => x"13070040",
         478 => x"b387e740",
         479 => x"6376f500",
         480 => x"13060500",
         481 => x"6ff05fd2",
         482 => x"ef109034",
         483 => x"9307c000",
         484 => x"2320f500",
         485 => x"1306f0ff",
         486 => x"6ff01fd1",
         487 => x"130e0500",
         488 => x"13830500",
         489 => x"13070000",
         490 => x"63dc0500",
         491 => x"b337a000",
         492 => x"3303b040",
         493 => x"3303f340",
         494 => x"330ea040",
         495 => x"1307f0ff",
         496 => x"63dc0600",
         497 => x"b337c000",
         498 => x"b306d040",
         499 => x"1347f7ff",
         500 => x"b386f640",
         501 => x"3306c040",
         502 => x"13080600",
         503 => x"93850600",
         504 => x"93080e00",
         505 => x"93070300",
         506 => x"63960622",
         507 => x"37450000",
         508 => x"1305c5a6",
         509 => x"6374c30e",
         510 => x"b7060100",
         511 => x"6376d60c",
         512 => x"93360610",
         513 => x"93b61600",
         514 => x"93963600",
         515 => x"b35ed600",
         516 => x"3305d501",
         517 => x"03450500",
         518 => x"b306d500",
         519 => x"13050002",
         520 => x"638ea600",
         521 => x"3305d540",
         522 => x"b317a300",
         523 => x"b356de00",
         524 => x"3318a600",
         525 => x"b3e7f600",
         526 => x"b318ae00",
         527 => x"13530801",
         528 => x"33d56702",
         529 => x"13160801",
         530 => x"13560601",
         531 => x"b3f76702",
         532 => x"330ea602",
         533 => x"93960701",
         534 => x"93d70801",
         535 => x"b3e7f600",
         536 => x"63fac701",
         537 => x"b307f800",
         538 => x"63f4c701",
         539 => x"63fa0719",
         540 => x"1305f5ff",
         541 => x"b387c741",
         542 => x"b3d66702",
         543 => x"93980801",
         544 => x"93d80801",
         545 => x"b3f76702",
         546 => x"3306d602",
         547 => x"93970701",
         548 => x"b3e8f800",
         549 => x"63fac800",
         550 => x"b3081801",
         551 => x"63f4c800",
         552 => x"63f60817",
         553 => x"9386f6ff",
         554 => x"13150501",
         555 => x"3365d500",
         556 => x"630a0700",
         557 => x"b337a000",
         558 => x"b305b040",
         559 => x"b385f540",
         560 => x"3305a040",
         561 => x"67800000",
         562 => x"b70e0001",
         563 => x"93068001",
         564 => x"e37ed6f3",
         565 => x"93060001",
         566 => x"6ff05ff3",
         567 => x"93060000",
         568 => x"630c0600",
         569 => x"b7070100",
         570 => x"637af604",
         571 => x"93360610",
         572 => x"93b61600",
         573 => x"93963600",
         574 => x"b357d600",
         575 => x"3305f500",
         576 => x"83470500",
         577 => x"93050002",
         578 => x"b387d700",
         579 => x"6392b704",
         580 => x"b307c340",
         581 => x"93051000",
         582 => x"13530801",
         583 => x"33d56702",
         584 => x"13160801",
         585 => x"13560601",
         586 => x"93d60801",
         587 => x"b3f76702",
         588 => x"330ea602",
         589 => x"93970701",
         590 => x"6ff05ff2",
         591 => x"b7070001",
         592 => x"93068001",
         593 => x"e37af6fa",
         594 => x"93060001",
         595 => x"6ff0dffa",
         596 => x"b385f540",
         597 => x"3318b600",
         598 => x"b356f300",
         599 => x"3313b300",
         600 => x"b357fe00",
         601 => x"b3e76700",
         602 => x"13530801",
         603 => x"b318be00",
         604 => x"b3d56602",
         605 => x"13150801",
         606 => x"13550501",
         607 => x"b3f66602",
         608 => x"330eb502",
         609 => x"13960601",
         610 => x"93d60701",
         611 => x"b3e6c600",
         612 => x"63fac601",
         613 => x"b306d800",
         614 => x"63f4c601",
         615 => x"63f60605",
         616 => x"9385f5ff",
         617 => x"b386c641",
         618 => x"33d66602",
         619 => x"93970701",
         620 => x"93d70701",
         621 => x"b3f66602",
         622 => x"3305c502",
         623 => x"93960601",
         624 => x"b3e7d700",
         625 => x"63faa700",
         626 => x"b307f800",
         627 => x"63f4a700",
         628 => x"63f20703",
         629 => x"1306f6ff",
         630 => x"93950501",
         631 => x"b387a740",
         632 => x"b3e5c500",
         633 => x"6ff05ff3",
         634 => x"9385e5ff",
         635 => x"b3860601",
         636 => x"6ff05ffb",
         637 => x"1306e6ff",
         638 => x"b3870701",
         639 => x"6ff0dffd",
         640 => x"1305e5ff",
         641 => x"b3870701",
         642 => x"6ff0dfe6",
         643 => x"9386e6ff",
         644 => x"6ff09fe9",
         645 => x"6364d318",
         646 => x"b7070100",
         647 => x"63f4f604",
         648 => x"93b50610",
         649 => x"93b51500",
         650 => x"93953500",
         651 => x"b7470000",
         652 => x"33d5b600",
         653 => x"9387c7a6",
         654 => x"b387a700",
         655 => x"83c70700",
         656 => x"930e0002",
         657 => x"b387b700",
         658 => x"6398d703",
         659 => x"3335ce00",
         660 => x"13351500",
         661 => x"b3b66600",
         662 => x"3365d500",
         663 => x"93050000",
         664 => x"6ff01fe5",
         665 => x"b7070001",
         666 => x"93058001",
         667 => x"e3f0f6fc",
         668 => x"93050001",
         669 => x"6ff09ffb",
         670 => x"b38efe40",
         671 => x"b355f600",
         672 => x"b396d601",
         673 => x"3358f300",
         674 => x"b3e6d500",
         675 => x"3313d301",
         676 => x"b357fe00",
         677 => x"b3e56700",
         678 => x"13d30601",
         679 => x"b3576802",
         680 => x"13950601",
         681 => x"13550501",
         682 => x"3316d601",
         683 => x"33786802",
         684 => x"330ff502",
         685 => x"93180801",
         686 => x"13d80501",
         687 => x"33681801",
         688 => x"637ae801",
         689 => x"33880601",
         690 => x"6374e801",
         691 => x"637cd80a",
         692 => x"9387f7ff",
         693 => x"3308e841",
         694 => x"b3586802",
         695 => x"93950501",
         696 => x"93d50501",
         697 => x"33786802",
         698 => x"33051503",
         699 => x"13180801",
         700 => x"b3e50501",
         701 => x"63faa500",
         702 => x"b385b600",
         703 => x"63f4a500",
         704 => x"63f8d508",
         705 => x"9388f8ff",
         706 => x"93970701",
         707 => x"13180601",
         708 => x"b385a540",
         709 => x"33e51701",
         710 => x"93980801",
         711 => x"93d80801",
         712 => x"93560501",
         713 => x"13580801",
         714 => x"13560601",
         715 => x"33830803",
         716 => x"33880603",
         717 => x"93570301",
         718 => x"b388c802",
         719 => x"b3880801",
         720 => x"b3871701",
         721 => x"b386c602",
         722 => x"63f60701",
         723 => x"37060100",
         724 => x"b386c600",
         725 => x"13d60701",
         726 => x"b306d600",
         727 => x"63e0d502",
         728 => x"13130301",
         729 => x"93970701",
         730 => x"13530301",
         731 => x"331ede01",
         732 => x"b3876700",
         733 => x"e374feee",
         734 => x"e392d5ee",
         735 => x"1305f5ff",
         736 => x"6ff0dfed",
         737 => x"9387e7ff",
         738 => x"3308d800",
         739 => x"6ff09ff4",
         740 => x"9388e8ff",
         741 => x"b385d500",
         742 => x"6ff01ff7",
         743 => x"93050000",
         744 => x"13050000",
         745 => x"6ff0dfd0",
         746 => x"13070600",
         747 => x"93880600",
         748 => x"13080500",
         749 => x"13830500",
         750 => x"63940624",
         751 => x"b7470000",
         752 => x"9387c7a6",
         753 => x"63f4c50e",
         754 => x"b7060100",
         755 => x"6370d60c",
         756 => x"93360610",
         757 => x"93b61600",
         758 => x"93963600",
         759 => x"335ed600",
         760 => x"b387c701",
         761 => x"83c70700",
         762 => x"b387d700",
         763 => x"93060002",
         764 => x"638ed700",
         765 => x"b386f640",
         766 => x"3393d500",
         767 => x"b357f500",
         768 => x"3317d600",
         769 => x"33e36700",
         770 => x"3318d500",
         771 => x"13550701",
         772 => x"b357a302",
         773 => x"93150701",
         774 => x"93d50501",
         775 => x"93560801",
         776 => x"3373a302",
         777 => x"3386f502",
         778 => x"13130301",
         779 => x"b3e66600",
         780 => x"63fac600",
         781 => x"b306d700",
         782 => x"63f4c600",
         783 => x"63f2e606",
         784 => x"9387f7ff",
         785 => x"b386c640",
         786 => x"33d6a602",
         787 => x"13180801",
         788 => x"13580801",
         789 => x"b3f6a602",
         790 => x"b385c502",
         791 => x"93960601",
         792 => x"3368d800",
         793 => x"637ab800",
         794 => x"33080701",
         795 => x"6374b800",
         796 => x"6374e818",
         797 => x"1306f6ff",
         798 => x"93970701",
         799 => x"b3e7c700",
         800 => x"13850700",
         801 => x"93850800",
         802 => x"67800000",
         803 => x"370e0001",
         804 => x"93068001",
         805 => x"e374c6f5",
         806 => x"93060001",
         807 => x"6ff01ff4",
         808 => x"9387e7ff",
         809 => x"b386e600",
         810 => x"6ff0dff9",
         811 => x"93060000",
         812 => x"630c0600",
         813 => x"b7060100",
         814 => x"6378d606",
         815 => x"93360610",
         816 => x"93b61600",
         817 => x"93963600",
         818 => x"b358d600",
         819 => x"b3871701",
         820 => x"83c70700",
         821 => x"b387d700",
         822 => x"93060002",
         823 => x"6390d706",
         824 => x"3386c540",
         825 => x"93081000",
         826 => x"13550701",
         827 => x"b357a602",
         828 => x"93150701",
         829 => x"93d50501",
         830 => x"93560801",
         831 => x"3376a602",
         832 => x"3383f502",
         833 => x"13160601",
         834 => x"b3e6c600",
         835 => x"63fa6600",
         836 => x"b306d700",
         837 => x"63f46600",
         838 => x"63fae60c",
         839 => x"9387f7ff",
         840 => x"b3866640",
         841 => x"6ff05ff2",
         842 => x"b7080001",
         843 => x"93068001",
         844 => x"e37c16f9",
         845 => x"93060001",
         846 => x"6ff01ff9",
         847 => x"3388f640",
         848 => x"33170601",
         849 => x"b3d6f500",
         850 => x"b3950501",
         851 => x"b357f500",
         852 => x"33180501",
         853 => x"13550701",
         854 => x"b3d8a602",
         855 => x"13160701",
         856 => x"13560601",
         857 => x"b3e7b700",
         858 => x"b3f6a602",
         859 => x"33031603",
         860 => x"93950601",
         861 => x"93d60701",
         862 => x"b3e6b600",
         863 => x"63fa6600",
         864 => x"b306d700",
         865 => x"63f46600",
         866 => x"63f6e604",
         867 => x"9388f8ff",
         868 => x"b3866640",
         869 => x"b3d5a602",
         870 => x"93970701",
         871 => x"93d70701",
         872 => x"b3f6a602",
         873 => x"3306b602",
         874 => x"93960601",
         875 => x"b3e7d700",
         876 => x"63fac700",
         877 => x"b307f700",
         878 => x"63f4c700",
         879 => x"63f2e702",
         880 => x"9385f5ff",
         881 => x"93980801",
         882 => x"3386c740",
         883 => x"b3e8b800",
         884 => x"6ff09ff1",
         885 => x"9388e8ff",
         886 => x"b386e600",
         887 => x"6ff05ffb",
         888 => x"9385e5ff",
         889 => x"b387e700",
         890 => x"6ff0dffd",
         891 => x"9387e7ff",
         892 => x"b386e600",
         893 => x"6ff0dff2",
         894 => x"1306e6ff",
         895 => x"6ff0dfe7",
         896 => x"63e4d518",
         897 => x"b7070100",
         898 => x"63f4f604",
         899 => x"93b70610",
         900 => x"93b71700",
         901 => x"93973700",
         902 => x"37470000",
         903 => x"33d8f600",
         904 => x"1307c7a6",
         905 => x"33070701",
         906 => x"03470700",
         907 => x"13080002",
         908 => x"3307f700",
         909 => x"63180703",
         910 => x"b337c500",
         911 => x"93b71700",
         912 => x"b3b6b600",
         913 => x"b3e7d700",
         914 => x"93080000",
         915 => x"6ff05fe3",
         916 => x"37070001",
         917 => x"93078001",
         918 => x"e3f0e6fc",
         919 => x"93070001",
         920 => x"6ff09ffb",
         921 => x"3308e840",
         922 => x"b358e600",
         923 => x"b3960601",
         924 => x"b3e8d800",
         925 => x"13de0801",
         926 => x"b3d6e500",
         927 => x"b3d7c603",
         928 => x"13930801",
         929 => x"13530301",
         930 => x"b3950501",
         931 => x"3357e500",
         932 => x"3367b700",
         933 => x"33160601",
         934 => x"b3f6c603",
         935 => x"b30ef302",
         936 => x"93950601",
         937 => x"93560701",
         938 => x"b3e6b600",
         939 => x"63fad601",
         940 => x"b386d800",
         941 => x"63f4d601",
         942 => x"63fc160b",
         943 => x"9387f7ff",
         944 => x"b386d641",
         945 => x"b3d5c603",
         946 => x"13170701",
         947 => x"13570701",
         948 => x"b3f6c603",
         949 => x"3303b302",
         950 => x"93960601",
         951 => x"3367d700",
         952 => x"637a6700",
         953 => x"3387e800",
         954 => x"63746700",
         955 => x"63781709",
         956 => x"9385f5ff",
         957 => x"93970701",
         958 => x"b3e7b700",
         959 => x"33076740",
         960 => x"93950501",
         961 => x"13130601",
         962 => x"93d50501",
         963 => x"93d80701",
         964 => x"13530301",
         965 => x"13560601",
         966 => x"338e6502",
         967 => x"33836802",
         968 => x"93560e01",
         969 => x"b385c502",
         970 => x"b3856500",
         971 => x"b386b600",
         972 => x"b388c802",
         973 => x"63f66600",
         974 => x"37060100",
         975 => x"b388c800",
         976 => x"13d60601",
         977 => x"33061601",
         978 => x"6360c702",
         979 => x"131e0e01",
         980 => x"93960601",
         981 => x"135e0e01",
         982 => x"33150501",
         983 => x"b386c601",
         984 => x"e374d5ee",
         985 => x"e312c7ee",
         986 => x"9387f7ff",
         987 => x"6ff0dfed",
         988 => x"9387e7ff",
         989 => x"b3861601",
         990 => x"6ff09ff4",
         991 => x"9385e5ff",
         992 => x"33071701",
         993 => x"6ff01ff7",
         994 => x"93080000",
         995 => x"93070000",
         996 => x"6ff01fcf",
         997 => x"13080600",
         998 => x"93070500",
         999 => x"13870500",
        1000 => x"63940624",
        1001 => x"b7460000",
        1002 => x"9386c6a6",
        1003 => x"63f8c50e",
        1004 => x"b7080100",
        1005 => x"637a160d",
        1006 => x"93380610",
        1007 => x"93b81800",
        1008 => x"93983800",
        1009 => x"33531601",
        1010 => x"b3866600",
        1011 => x"83c60600",
        1012 => x"13030002",
        1013 => x"b3861601",
        1014 => x"b308d340",
        1015 => x"638c6600",
        1016 => x"33971501",
        1017 => x"b356d500",
        1018 => x"33181601",
        1019 => x"33e7e600",
        1020 => x"b3171501",
        1021 => x"13550801",
        1022 => x"b356a702",
        1023 => x"13130801",
        1024 => x"13530301",
        1025 => x"3377a702",
        1026 => x"b3866602",
        1027 => x"93150701",
        1028 => x"13d70701",
        1029 => x"3367b700",
        1030 => x"6370d702",
        1031 => x"3307e800",
        1032 => x"b3350701",
        1033 => x"3336d700",
        1034 => x"93b51500",
        1035 => x"3376b600",
        1036 => x"33060603",
        1037 => x"3307e600",
        1038 => x"3307d740",
        1039 => x"b356a702",
        1040 => x"3377a702",
        1041 => x"b3866602",
        1042 => x"13950701",
        1043 => x"13170701",
        1044 => x"13550501",
        1045 => x"3365e500",
        1046 => x"6370d502",
        1047 => x"3305a800",
        1048 => x"33370501",
        1049 => x"b337d500",
        1050 => x"13371700",
        1051 => x"b3f7e700",
        1052 => x"b3870703",
        1053 => x"3385a700",
        1054 => x"3305d540",
        1055 => x"33551501",
        1056 => x"93050000",
        1057 => x"67800000",
        1058 => x"37030001",
        1059 => x"93088001",
        1060 => x"e37a66f2",
        1061 => x"93080001",
        1062 => x"6ff0dff2",
        1063 => x"13070000",
        1064 => x"630c0600",
        1065 => x"37070100",
        1066 => x"6374e608",
        1067 => x"13370610",
        1068 => x"13371700",
        1069 => x"13173700",
        1070 => x"b358e600",
        1071 => x"b3861601",
        1072 => x"83c60600",
        1073 => x"b386e600",
        1074 => x"13070002",
        1075 => x"b308d740",
        1076 => x"639ae606",
        1077 => x"b386c540",
        1078 => x"93550801",
        1079 => x"33d6b602",
        1080 => x"13130801",
        1081 => x"13530301",
        1082 => x"13d70701",
        1083 => x"b3f6b602",
        1084 => x"33066602",
        1085 => x"93960601",
        1086 => x"3367d700",
        1087 => x"6370c702",
        1088 => x"3307e800",
        1089 => x"33350701",
        1090 => x"b336c700",
        1091 => x"13351500",
        1092 => x"b3f6a600",
        1093 => x"b3860603",
        1094 => x"3387e600",
        1095 => x"3307c740",
        1096 => x"b356b702",
        1097 => x"3377b702",
        1098 => x"b3866602",
        1099 => x"6ff0dff1",
        1100 => x"b7080001",
        1101 => x"13078001",
        1102 => x"e37016f9",
        1103 => x"13070001",
        1104 => x"6ff09ff7",
        1105 => x"33181601",
        1106 => x"33d7d500",
        1107 => x"b3171501",
        1108 => x"b3951501",
        1109 => x"b356d500",
        1110 => x"13550801",
        1111 => x"b3e6b600",
        1112 => x"b355a702",
        1113 => x"131e0801",
        1114 => x"135e0e01",
        1115 => x"3377a702",
        1116 => x"b385c503",
        1117 => x"13160701",
        1118 => x"13d70601",
        1119 => x"3367c700",
        1120 => x"6370b702",
        1121 => x"3307e800",
        1122 => x"33330701",
        1123 => x"3336b700",
        1124 => x"13331300",
        1125 => x"33766600",
        1126 => x"33060603",
        1127 => x"3307e600",
        1128 => x"3307b740",
        1129 => x"3356a702",
        1130 => x"93960601",
        1131 => x"93d60601",
        1132 => x"3377a702",
        1133 => x"3306c603",
        1134 => x"13170701",
        1135 => x"b3e6e600",
        1136 => x"63f0c602",
        1137 => x"b306d800",
        1138 => x"b3b50601",
        1139 => x"33b7c600",
        1140 => x"93b51500",
        1141 => x"3377b700",
        1142 => x"33070703",
        1143 => x"b306d700",
        1144 => x"b386c640",
        1145 => x"6ff05fef",
        1146 => x"63e6d51a",
        1147 => x"37080100",
        1148 => x"63fc0605",
        1149 => x"93b80610",
        1150 => x"93b81800",
        1151 => x"93983800",
        1152 => x"37480000",
        1153 => x"33d31601",
        1154 => x"1308c8a6",
        1155 => x"33086800",
        1156 => x"03480800",
        1157 => x"33081801",
        1158 => x"93080002",
        1159 => x"63101805",
        1160 => x"6374c500",
        1161 => x"63fcb600",
        1162 => x"3307c540",
        1163 => x"93070700",
        1164 => x"b386d540",
        1165 => x"3337e500",
        1166 => x"3387e640",
        1167 => x"13850700",
        1168 => x"93050700",
        1169 => x"67800000",
        1170 => x"37080001",
        1171 => x"93088001",
        1172 => x"e3f806fb",
        1173 => x"93080001",
        1174 => x"6ff09ffa",
        1175 => x"b3880841",
        1176 => x"b3961601",
        1177 => x"33530601",
        1178 => x"3363d300",
        1179 => x"33d70501",
        1180 => x"935e0301",
        1181 => x"b356d703",
        1182 => x"131e0301",
        1183 => x"135e0e01",
        1184 => x"b3971501",
        1185 => x"b3550501",
        1186 => x"b3e5f500",
        1187 => x"93d70501",
        1188 => x"33161601",
        1189 => x"33151501",
        1190 => x"3377d703",
        1191 => x"330fde02",
        1192 => x"13170701",
        1193 => x"b3e7e700",
        1194 => x"63fae701",
        1195 => x"b307f300",
        1196 => x"63f4e701",
        1197 => x"63f2670e",
        1198 => x"9386f6ff",
        1199 => x"b387e741",
        1200 => x"33d7d703",
        1201 => x"93950501",
        1202 => x"93d50501",
        1203 => x"b3f7d703",
        1204 => x"330eee02",
        1205 => x"93970701",
        1206 => x"b3e5f500",
        1207 => x"63fac501",
        1208 => x"b305b300",
        1209 => x"63f4c501",
        1210 => x"63fe650a",
        1211 => x"1307f7ff",
        1212 => x"93960601",
        1213 => x"b3e6e600",
        1214 => x"b385c541",
        1215 => x"13170701",
        1216 => x"131e0601",
        1217 => x"93570601",
        1218 => x"13570701",
        1219 => x"93d60601",
        1220 => x"135e0e01",
        1221 => x"b30ec703",
        1222 => x"338ec603",
        1223 => x"3307f702",
        1224 => x"b386f602",
        1225 => x"b307c701",
        1226 => x"13d70e01",
        1227 => x"3307f700",
        1228 => x"6376c701",
        1229 => x"b7070100",
        1230 => x"b386f600",
        1231 => x"93570701",
        1232 => x"939e0e01",
        1233 => x"13170701",
        1234 => x"93de0e01",
        1235 => x"b387d700",
        1236 => x"3307d701",
        1237 => x"63e6f500",
        1238 => x"637ee500",
        1239 => x"639cf500",
        1240 => x"3306c740",
        1241 => x"b336c700",
        1242 => x"b3866600",
        1243 => x"13070600",
        1244 => x"b387d740",
        1245 => x"3307e540",
        1246 => x"3335e500",
        1247 => x"b385f540",
        1248 => x"b385a540",
        1249 => x"33980501",
        1250 => x"33571701",
        1251 => x"3365e800",
        1252 => x"b3d51501",
        1253 => x"67800000",
        1254 => x"9386e6ff",
        1255 => x"b3876700",
        1256 => x"6ff0dff1",
        1257 => x"1307e7ff",
        1258 => x"b3856500",
        1259 => x"6ff05ff4",
        1260 => x"13030500",
        1261 => x"630a0600",
        1262 => x"2300b300",
        1263 => x"1306f6ff",
        1264 => x"13031300",
        1265 => x"e31a06fe",
        1266 => x"67800000",
        1267 => x"13030500",
        1268 => x"630e0600",
        1269 => x"83830500",
        1270 => x"23007300",
        1271 => x"1306f6ff",
        1272 => x"13031300",
        1273 => x"93851500",
        1274 => x"e31606fe",
        1275 => x"67800000",
        1276 => x"630c0602",
        1277 => x"13030500",
        1278 => x"93061000",
        1279 => x"636ab500",
        1280 => x"9306f0ff",
        1281 => x"1307f6ff",
        1282 => x"3303e300",
        1283 => x"b385e500",
        1284 => x"83830500",
        1285 => x"23007300",
        1286 => x"1306f6ff",
        1287 => x"3303d300",
        1288 => x"b385d500",
        1289 => x"e31606fe",
        1290 => x"67800000",
        1291 => x"370700f0",
        1292 => x"13070710",
        1293 => x"83274700",
        1294 => x"93f78700",
        1295 => x"e38c07fe",
        1296 => x"03258700",
        1297 => x"1375f50f",
        1298 => x"67800000",
        1299 => x"f32710fc",
        1300 => x"63960700",
        1301 => x"b7f7fa02",
        1302 => x"93870708",
        1303 => x"63060500",
        1304 => x"33d5a702",
        1305 => x"1305f5ff",
        1306 => x"b70700f0",
        1307 => x"23a6a710",
        1308 => x"23a0b710",
        1309 => x"23a20710",
        1310 => x"67800000",
        1311 => x"370700f0",
        1312 => x"1375f50f",
        1313 => x"13070710",
        1314 => x"2324a700",
        1315 => x"83274700",
        1316 => x"93f70701",
        1317 => x"e38c07fe",
        1318 => x"67800000",
        1319 => x"630e0502",
        1320 => x"130101ff",
        1321 => x"23248100",
        1322 => x"23261100",
        1323 => x"13040500",
        1324 => x"03450500",
        1325 => x"630a0500",
        1326 => x"13041400",
        1327 => x"eff01ffc",
        1328 => x"03450400",
        1329 => x"e31a05fe",
        1330 => x"8320c100",
        1331 => x"03248100",
        1332 => x"13010101",
        1333 => x"67800000",
        1334 => x"67800000",
        1335 => x"130101fd",
        1336 => x"23261102",
        1337 => x"232a0100",
        1338 => x"232c0100",
        1339 => x"232e0100",
        1340 => x"63000508",
        1341 => x"93070500",
        1342 => x"63400506",
        1343 => x"b7d5cccc",
        1344 => x"13850700",
        1345 => x"9385d5cc",
        1346 => x"93064101",
        1347 => x"93089000",
        1348 => x"b337b502",
        1349 => x"13060500",
        1350 => x"13880600",
        1351 => x"9386f6ff",
        1352 => x"93d73700",
        1353 => x"13972700",
        1354 => x"3307f700",
        1355 => x"13171700",
        1356 => x"3305e540",
        1357 => x"13050503",
        1358 => x"a385a600",
        1359 => x"13850700",
        1360 => x"e3e8c8fc",
        1361 => x"1305a800",
        1362 => x"eff05ff5",
        1363 => x"8320c102",
        1364 => x"13010103",
        1365 => x"67800000",
        1366 => x"2326a100",
        1367 => x"1305d002",
        1368 => x"eff0dff1",
        1369 => x"8327c100",
        1370 => x"b307f040",
        1371 => x"6ff01ff9",
        1372 => x"13050003",
        1373 => x"eff09ff0",
        1374 => x"8320c102",
        1375 => x"13010103",
        1376 => x"67800000",
        1377 => x"130101ff",
        1378 => x"23261100",
        1379 => x"23248100",
        1380 => x"732430f1",
        1381 => x"1355c401",
        1382 => x"63140508",
        1383 => x"13558401",
        1384 => x"1375f500",
        1385 => x"13050503",
        1386 => x"eff05fed",
        1387 => x"1305e002",
        1388 => x"eff0dfec",
        1389 => x"13554401",
        1390 => x"1375f500",
        1391 => x"631e0508",
        1392 => x"13550401",
        1393 => x"1375f500",
        1394 => x"13050503",
        1395 => x"eff01feb",
        1396 => x"1305e002",
        1397 => x"eff09fea",
        1398 => x"1355c400",
        1399 => x"1375f500",
        1400 => x"63160506",
        1401 => x"13558400",
        1402 => x"1375f500",
        1403 => x"13050503",
        1404 => x"eff0dfe8",
        1405 => x"1305e002",
        1406 => x"eff05fe8",
        1407 => x"13554400",
        1408 => x"1375f500",
        1409 => x"63140502",
        1410 => x"1375f400",
        1411 => x"03248100",
        1412 => x"8320c100",
        1413 => x"13050503",
        1414 => x"13010101",
        1415 => x"6ff01fe6",
        1416 => x"13050503",
        1417 => x"eff09fe5",
        1418 => x"6ff05ff7",
        1419 => x"13050503",
        1420 => x"eff0dfe4",
        1421 => x"1375f400",
        1422 => x"03248100",
        1423 => x"8320c100",
        1424 => x"13050503",
        1425 => x"13010101",
        1426 => x"6ff05fe3",
        1427 => x"13050503",
        1428 => x"eff0dfe2",
        1429 => x"6ff01ff9",
        1430 => x"13050503",
        1431 => x"eff01fe2",
        1432 => x"6ff01ff6",
        1433 => x"130101f9",
        1434 => x"23229106",
        1435 => x"23202107",
        1436 => x"23261106",
        1437 => x"23248106",
        1438 => x"232e3105",
        1439 => x"232a5105",
        1440 => x"23286105",
        1441 => x"23267105",
        1442 => x"23248105",
        1443 => x"23229105",
        1444 => x"2320a105",
        1445 => x"13890500",
        1446 => x"93040500",
        1447 => x"f32a00fc",
        1448 => x"b7070008",
        1449 => x"232c0100",
        1450 => x"232e0100",
        1451 => x"23200102",
        1452 => x"23220102",
        1453 => x"23240102",
        1454 => x"23260102",
        1455 => x"23280102",
        1456 => x"232a0102",
        1457 => x"232c0102",
        1458 => x"232e0102",
        1459 => x"b3fafa00",
        1460 => x"732410fc",
        1461 => x"63160400",
        1462 => x"37f4fa02",
        1463 => x"13040408",
        1464 => x"97f2ffff",
        1465 => x"938242c2",
        1466 => x"73905230",
        1467 => x"37c50100",
        1468 => x"13050520",
        1469 => x"93059000",
        1470 => x"eff05fd5",
        1471 => x"b716b7d1",
        1472 => x"93869675",
        1473 => x"b336d402",
        1474 => x"37353e05",
        1475 => x"13576400",
        1476 => x"130535d6",
        1477 => x"b727d96f",
        1478 => x"938757d8",
        1479 => x"13561400",
        1480 => x"b70500f0",
        1481 => x"1306f6ff",
        1482 => x"23a6c560",
        1483 => x"3337a702",
        1484 => x"93d6d600",
        1485 => x"13051001",
        1486 => x"23a0a560",
        1487 => x"9386f6ff",
        1488 => x"23a8d570",
        1489 => x"b7260000",
        1490 => x"9386f670",
        1491 => x"23a6d570",
        1492 => x"13860500",
        1493 => x"b337f402",
        1494 => x"13576700",
        1495 => x"1307f7ff",
        1496 => x"23a0a570",
        1497 => x"13170701",
        1498 => x"93058070",
        1499 => x"2320b640",
        1500 => x"13678700",
        1501 => x"2320e620",
        1502 => x"1307a007",
        1503 => x"93d73701",
        1504 => x"9387f7ff",
        1505 => x"93970701",
        1506 => x"93e7c700",
        1507 => x"2320f630",
        1508 => x"232ce600",
        1509 => x"f3224030",
        1510 => x"93e20208",
        1511 => x"73904230",
        1512 => x"f3224030",
        1513 => x"93e28200",
        1514 => x"73904230",
        1515 => x"b7220000",
        1516 => x"93828280",
        1517 => x"73900230",
        1518 => x"b7490000",
        1519 => x"1385c9b8",
        1520 => x"eff0dfcd",
        1521 => x"635a9002",
        1522 => x"232c4105",
        1523 => x"9384f4ff",
        1524 => x"9389c9b8",
        1525 => x"130af0ff",
        1526 => x"03250900",
        1527 => x"9384f4ff",
        1528 => x"13094900",
        1529 => x"eff09fcb",
        1530 => x"13850900",
        1531 => x"eff01fcb",
        1532 => x"e39444ff",
        1533 => x"032a8105",
        1534 => x"37450000",
        1535 => x"130505b9",
        1536 => x"eff0dfc9",
        1537 => x"13050400",
        1538 => x"eff05fcd",
        1539 => x"37450000",
        1540 => x"130545ba",
        1541 => x"eff09fc8",
        1542 => x"eff0dfd6",
        1543 => x"37450000",
        1544 => x"1305c5bb",
        1545 => x"eff09fc7",
        1546 => x"63980a22",
        1547 => x"b7040010",
        1548 => x"37f4eeee",
        1549 => x"b7998888",
        1550 => x"9384f4ff",
        1551 => x"93899988",
        1552 => x"1304f4ee",
        1553 => x"374b0000",
        1554 => x"371c0000",
        1555 => x"37f9eeee",
        1556 => x"130c0c2c",
        1557 => x"1309e9ee",
        1558 => x"6f00c000",
        1559 => x"130cfcff",
        1560 => x"63040c1a",
        1561 => x"93050000",
        1562 => x"13058100",
        1563 => x"ef001030",
        1564 => x"e31605fe",
        1565 => x"832c8100",
        1566 => x"8325c100",
        1567 => x"37160000",
        1568 => x"93d7cc01",
        1569 => x"13974500",
        1570 => x"b307f700",
        1571 => x"33f79700",
        1572 => x"b3f79c00",
        1573 => x"b387e700",
        1574 => x"13d78501",
        1575 => x"b387e700",
        1576 => x"13d7f541",
        1577 => x"1375d700",
        1578 => x"b387a700",
        1579 => x"33b83703",
        1580 => x"137727ff",
        1581 => x"130606e1",
        1582 => x"93060000",
        1583 => x"13850c00",
        1584 => x"130cfcff",
        1585 => x"13583800",
        1586 => x"93184800",
        1587 => x"33880841",
        1588 => x"b3870741",
        1589 => x"b387e700",
        1590 => x"13d7f741",
        1591 => x"b387fc40",
        1592 => x"33b8fc00",
        1593 => x"3387e540",
        1594 => x"33070741",
        1595 => x"33078702",
        1596 => x"33882703",
        1597 => x"33070701",
        1598 => x"33b88702",
        1599 => x"b3878702",
        1600 => x"33070701",
        1601 => x"1358f741",
        1602 => x"13783800",
        1603 => x"b307f800",
        1604 => x"33b80701",
        1605 => x"3308e800",
        1606 => x"1317e801",
        1607 => x"93d72700",
        1608 => x"b307f700",
        1609 => x"93582840",
        1610 => x"13d7c701",
        1611 => x"13934800",
        1612 => x"3307e300",
        1613 => x"33739700",
        1614 => x"33f79700",
        1615 => x"33076700",
        1616 => x"1358f841",
        1617 => x"13d38801",
        1618 => x"33076700",
        1619 => x"1373d800",
        1620 => x"33076700",
        1621 => x"33333703",
        1622 => x"137828ff",
        1623 => x"939b4700",
        1624 => x"b38bfb40",
        1625 => x"939b2b00",
        1626 => x"13533300",
        1627 => x"131e4300",
        1628 => x"33036e40",
        1629 => x"33076740",
        1630 => x"33070701",
        1631 => x"1358f741",
        1632 => x"3387e740",
        1633 => x"33880841",
        1634 => x"b3b8e700",
        1635 => x"33081841",
        1636 => x"33032703",
        1637 => x"33088802",
        1638 => x"b3388702",
        1639 => x"33086800",
        1640 => x"33078702",
        1641 => x"33081801",
        1642 => x"9358f841",
        1643 => x"93f83800",
        1644 => x"3387e800",
        1645 => x"b3381701",
        1646 => x"b3880801",
        1647 => x"9398e801",
        1648 => x"13572700",
        1649 => x"3387e800",
        1650 => x"13184700",
        1651 => x"3307e840",
        1652 => x"13172700",
        1653 => x"338de740",
        1654 => x"efe05fdc",
        1655 => x"83260101",
        1656 => x"13070500",
        1657 => x"33887c41",
        1658 => x"93070d00",
        1659 => x"13860c00",
        1660 => x"93054bc2",
        1661 => x"13058101",
        1662 => x"ef008047",
        1663 => x"13058101",
        1664 => x"eff0dfa9",
        1665 => x"e3100ce6",
        1666 => x"63940a00",
        1667 => x"73001000",
        1668 => x"b70700f0",
        1669 => x"1307f00f",
        1670 => x"23a4e740",
        1671 => x"370700f0",
        1672 => x"83260720",
        1673 => x"13060009",
        1674 => x"93070700",
        1675 => x"93e60630",
        1676 => x"2320d720",
        1677 => x"2324c720",
        1678 => x"83260730",
        1679 => x"371700f0",
        1680 => x"93e60630",
        1681 => x"23a0d730",
        1682 => x"23a4c730",
        1683 => x"93071000",
        1684 => x"2320f790",
        1685 => x"6ff05fdf",
        1686 => x"37450000",
        1687 => x"1305c5be",
        1688 => x"eff0dfa3",
        1689 => x"6ff09fdc",
        1690 => x"130101ff",
        1691 => x"23248100",
        1692 => x"23261100",
        1693 => x"93070000",
        1694 => x"13040500",
        1695 => x"63880700",
        1696 => x"93050000",
        1697 => x"97000000",
        1698 => x"e7000000",
        1699 => x"83a74187",
        1700 => x"63840700",
        1701 => x"e7800700",
        1702 => x"13050400",
        1703 => x"ef101044",
        1704 => x"13050000",
        1705 => x"67800000",
        1706 => x"130101ff",
        1707 => x"23248100",
        1708 => x"23261100",
        1709 => x"13040500",
        1710 => x"2316b500",
        1711 => x"2317c500",
        1712 => x"23200500",
        1713 => x"23220500",
        1714 => x"23240500",
        1715 => x"23220506",
        1716 => x"23280500",
        1717 => x"232a0500",
        1718 => x"232c0500",
        1719 => x"13068000",
        1720 => x"93050000",
        1721 => x"1305c505",
        1722 => x"eff09f8c",
        1723 => x"b7270000",
        1724 => x"938747ee",
        1725 => x"2322f402",
        1726 => x"b7270000",
        1727 => x"9387c7f3",
        1728 => x"2324f402",
        1729 => x"b7270000",
        1730 => x"938707fc",
        1731 => x"2326f402",
        1732 => x"b7270000",
        1733 => x"93878701",
        1734 => x"8320c100",
        1735 => x"23208402",
        1736 => x"2328f402",
        1737 => x"03248100",
        1738 => x"13010101",
        1739 => x"67800000",
        1740 => x"b7350000",
        1741 => x"37050020",
        1742 => x"13868181",
        1743 => x"9385c547",
        1744 => x"13054502",
        1745 => x"6f00c021",
        1746 => x"83254500",
        1747 => x"130101ff",
        1748 => x"b7070020",
        1749 => x"23248100",
        1750 => x"23261100",
        1751 => x"93878708",
        1752 => x"13040500",
        1753 => x"6384f500",
        1754 => x"ef105011",
        1755 => x"83258400",
        1756 => x"9387018f",
        1757 => x"6386f500",
        1758 => x"13050400",
        1759 => x"ef101010",
        1760 => x"8325c400",
        1761 => x"93878195",
        1762 => x"638cf500",
        1763 => x"13050400",
        1764 => x"03248100",
        1765 => x"8320c100",
        1766 => x"13010101",
        1767 => x"6f10100e",
        1768 => x"8320c100",
        1769 => x"03248100",
        1770 => x"13010101",
        1771 => x"67800000",
        1772 => x"b7270000",
        1773 => x"37050020",
        1774 => x"130101ff",
        1775 => x"938707b3",
        1776 => x"13060000",
        1777 => x"93054000",
        1778 => x"13058508",
        1779 => x"23261100",
        1780 => x"23aaf186",
        1781 => x"eff05fed",
        1782 => x"13061000",
        1783 => x"93059000",
        1784 => x"1385018f",
        1785 => x"eff05fec",
        1786 => x"8320c100",
        1787 => x"13062000",
        1788 => x"93052001",
        1789 => x"13858195",
        1790 => x"13010101",
        1791 => x"6ff0dfea",
        1792 => x"13050000",
        1793 => x"67800000",
        1794 => x"83a74187",
        1795 => x"130101ff",
        1796 => x"23202101",
        1797 => x"23261100",
        1798 => x"23248100",
        1799 => x"23229100",
        1800 => x"13090500",
        1801 => x"63940700",
        1802 => x"eff09ff8",
        1803 => x"93848181",
        1804 => x"03a48400",
        1805 => x"83a74400",
        1806 => x"9387f7ff",
        1807 => x"63d80702",
        1808 => x"03a40400",
        1809 => x"6310040c",
        1810 => x"9305c01a",
        1811 => x"13050900",
        1812 => x"ef00900a",
        1813 => x"13040500",
        1814 => x"63140508",
        1815 => x"23a00400",
        1816 => x"9307c000",
        1817 => x"2320f900",
        1818 => x"6f004005",
        1819 => x"0317c400",
        1820 => x"63140706",
        1821 => x"b707ffff",
        1822 => x"93871700",
        1823 => x"23220406",
        1824 => x"23200400",
        1825 => x"23220400",
        1826 => x"23240400",
        1827 => x"2326f400",
        1828 => x"23280400",
        1829 => x"232a0400",
        1830 => x"232c0400",
        1831 => x"13068000",
        1832 => x"93050000",
        1833 => x"1305c405",
        1834 => x"eff08ff0",
        1835 => x"232a0402",
        1836 => x"232c0402",
        1837 => x"23240404",
        1838 => x"23260404",
        1839 => x"8320c100",
        1840 => x"13050400",
        1841 => x"03248100",
        1842 => x"83244100",
        1843 => x"03290100",
        1844 => x"13010101",
        1845 => x"67800000",
        1846 => x"13048406",
        1847 => x"6ff0dff5",
        1848 => x"93074000",
        1849 => x"23200500",
        1850 => x"2322f500",
        1851 => x"1305c500",
        1852 => x"2324a400",
        1853 => x"1306001a",
        1854 => x"93050000",
        1855 => x"eff04feb",
        1856 => x"23a08400",
        1857 => x"93040400",
        1858 => x"6ff09ff2",
        1859 => x"83270502",
        1860 => x"639e0700",
        1861 => x"b7270000",
        1862 => x"938787b4",
        1863 => x"2320f502",
        1864 => x"83a74187",
        1865 => x"63940700",
        1866 => x"6ff09fe8",
        1867 => x"67800000",
        1868 => x"67800000",
        1869 => x"67800000",
        1870 => x"b7250000",
        1871 => x"13868181",
        1872 => x"938505aa",
        1873 => x"13050000",
        1874 => x"6f008001",
        1875 => x"b7250000",
        1876 => x"13868181",
        1877 => x"938505c0",
        1878 => x"13050000",
        1879 => x"6f004000",
        1880 => x"130101fd",
        1881 => x"23248102",
        1882 => x"23202103",
        1883 => x"232e3101",
        1884 => x"232c4101",
        1885 => x"232a5101",
        1886 => x"23261102",
        1887 => x"23229102",
        1888 => x"130a0500",
        1889 => x"938a0500",
        1890 => x"13040000",
        1891 => x"13091000",
        1892 => x"9309f0ff",
        1893 => x"83258600",
        1894 => x"83244600",
        1895 => x"9384f4ff",
        1896 => x"63da0402",
        1897 => x"03260600",
        1898 => x"e31606fe",
        1899 => x"8320c102",
        1900 => x"13050400",
        1901 => x"03248102",
        1902 => x"83244102",
        1903 => x"03290102",
        1904 => x"8329c101",
        1905 => x"032a8101",
        1906 => x"832a4101",
        1907 => x"13010103",
        1908 => x"67800000",
        1909 => x"83d7c500",
        1910 => x"6374f902",
        1911 => x"8397e500",
        1912 => x"63803703",
        1913 => x"13050a00",
        1914 => x"2326c100",
        1915 => x"2324b100",
        1916 => x"e7800a00",
        1917 => x"0326c100",
        1918 => x"83258100",
        1919 => x"3364a400",
        1920 => x"93858506",
        1921 => x"6ff09ff9",
        1922 => x"130101f6",
        1923 => x"232af108",
        1924 => x"b7070080",
        1925 => x"9387f7ff",
        1926 => x"232ef100",
        1927 => x"2328f100",
        1928 => x"b707ffff",
        1929 => x"2326d108",
        1930 => x"2324b100",
        1931 => x"232cb100",
        1932 => x"93878720",
        1933 => x"9306c108",
        1934 => x"93058100",
        1935 => x"232e1106",
        1936 => x"232af100",
        1937 => x"2328e108",
        1938 => x"232c0109",
        1939 => x"232e1109",
        1940 => x"23260106",
        1941 => x"2322d100",
        1942 => x"ef00103a",
        1943 => x"83278100",
        1944 => x"23800700",
        1945 => x"8320c107",
        1946 => x"1301010a",
        1947 => x"67800000",
        1948 => x"130101f6",
        1949 => x"232af108",
        1950 => x"b7070080",
        1951 => x"9387f7ff",
        1952 => x"232ef100",
        1953 => x"2328f100",
        1954 => x"b707ffff",
        1955 => x"93878720",
        1956 => x"232af100",
        1957 => x"2324a100",
        1958 => x"232ca100",
        1959 => x"03a50187",
        1960 => x"2324c108",
        1961 => x"2326d108",
        1962 => x"13860500",
        1963 => x"93068108",
        1964 => x"93058100",
        1965 => x"232e1106",
        1966 => x"2328e108",
        1967 => x"232c0109",
        1968 => x"232e1109",
        1969 => x"23260106",
        1970 => x"2322d100",
        1971 => x"ef00d032",
        1972 => x"83278100",
        1973 => x"23800700",
        1974 => x"8320c107",
        1975 => x"1301010a",
        1976 => x"67800000",
        1977 => x"130101ff",
        1978 => x"23248100",
        1979 => x"13840500",
        1980 => x"8395e500",
        1981 => x"23261100",
        1982 => x"ef008033",
        1983 => x"63400502",
        1984 => x"83274405",
        1985 => x"b387a700",
        1986 => x"232af404",
        1987 => x"8320c100",
        1988 => x"03248100",
        1989 => x"13010101",
        1990 => x"67800000",
        1991 => x"8357c400",
        1992 => x"37f7ffff",
        1993 => x"1307f7ff",
        1994 => x"b3f7e700",
        1995 => x"2316f400",
        1996 => x"6ff0dffd",
        1997 => x"13050000",
        1998 => x"67800000",
        1999 => x"83d7c500",
        2000 => x"130101fe",
        2001 => x"232c8100",
        2002 => x"232a9100",
        2003 => x"23282101",
        2004 => x"23263101",
        2005 => x"232e1100",
        2006 => x"93f70710",
        2007 => x"93040500",
        2008 => x"13840500",
        2009 => x"13090600",
        2010 => x"93890600",
        2011 => x"638a0700",
        2012 => x"8395e500",
        2013 => x"93062000",
        2014 => x"13060000",
        2015 => x"ef004026",
        2016 => x"8357c400",
        2017 => x"37f7ffff",
        2018 => x"1307f7ff",
        2019 => x"b3f7e700",
        2020 => x"8315e400",
        2021 => x"2316f400",
        2022 => x"03248101",
        2023 => x"8320c101",
        2024 => x"93860900",
        2025 => x"13060900",
        2026 => x"8329c100",
        2027 => x"03290101",
        2028 => x"13850400",
        2029 => x"83244101",
        2030 => x"13010102",
        2031 => x"6f00402c",
        2032 => x"130101ff",
        2033 => x"23248100",
        2034 => x"13840500",
        2035 => x"8395e500",
        2036 => x"23261100",
        2037 => x"ef00c020",
        2038 => x"1307f0ff",
        2039 => x"8317c400",
        2040 => x"6312e502",
        2041 => x"13070580",
        2042 => x"13070780",
        2043 => x"b3f7e700",
        2044 => x"2316f400",
        2045 => x"8320c100",
        2046 => x"03248100",
        2047 => x"13010101",
        2048 => x"67800000",
        2049 => x"37170000",
        2050 => x"b3e7e700",
        2051 => x"2316f400",
        2052 => x"232aa404",
        2053 => x"6ff01ffe",
        2054 => x"8395e500",
        2055 => x"6f004000",
        2056 => x"130101ff",
        2057 => x"23248100",
        2058 => x"23229100",
        2059 => x"93040500",
        2060 => x"13850500",
        2061 => x"23261100",
        2062 => x"23ac0186",
        2063 => x"ef100066",
        2064 => x"9307f0ff",
        2065 => x"6318f500",
        2066 => x"83a78187",
        2067 => x"63840700",
        2068 => x"23a0f400",
        2069 => x"8320c100",
        2070 => x"03248100",
        2071 => x"83244100",
        2072 => x"13010101",
        2073 => x"67800000",
        2074 => x"83a70187",
        2075 => x"6388a716",
        2076 => x"8327c501",
        2077 => x"130101fe",
        2078 => x"232c8100",
        2079 => x"232e1100",
        2080 => x"232a9100",
        2081 => x"23282101",
        2082 => x"23263101",
        2083 => x"13040500",
        2084 => x"63840708",
        2085 => x"83a7c700",
        2086 => x"638c0702",
        2087 => x"93040000",
        2088 => x"13090008",
        2089 => x"8327c401",
        2090 => x"83a7c700",
        2091 => x"b3879700",
        2092 => x"83a50700",
        2093 => x"63980504",
        2094 => x"93844400",
        2095 => x"e39424ff",
        2096 => x"8327c401",
        2097 => x"13050400",
        2098 => x"83a5c700",
        2099 => x"ef00002b",
        2100 => x"8327c401",
        2101 => x"83a50700",
        2102 => x"63860500",
        2103 => x"13050400",
        2104 => x"ef00c029",
        2105 => x"8327c401",
        2106 => x"83a48700",
        2107 => x"63860402",
        2108 => x"93850400",
        2109 => x"13050400",
        2110 => x"83a40400",
        2111 => x"ef000028",
        2112 => x"6ff0dffe",
        2113 => x"83a90500",
        2114 => x"13050400",
        2115 => x"ef000027",
        2116 => x"93850900",
        2117 => x"6ff01ffa",
        2118 => x"83254401",
        2119 => x"63860500",
        2120 => x"13050400",
        2121 => x"ef008025",
        2122 => x"8325c401",
        2123 => x"63860500",
        2124 => x"13050400",
        2125 => x"ef008024",
        2126 => x"83250403",
        2127 => x"63860500",
        2128 => x"13050400",
        2129 => x"ef008023",
        2130 => x"83254403",
        2131 => x"63860500",
        2132 => x"13050400",
        2133 => x"ef008022",
        2134 => x"83258403",
        2135 => x"63860500",
        2136 => x"13050400",
        2137 => x"ef008021",
        2138 => x"83258404",
        2139 => x"63860500",
        2140 => x"13050400",
        2141 => x"ef008020",
        2142 => x"83254404",
        2143 => x"63860500",
        2144 => x"13050400",
        2145 => x"ef00801f",
        2146 => x"8325c402",
        2147 => x"63860500",
        2148 => x"13050400",
        2149 => x"ef00801e",
        2150 => x"83270402",
        2151 => x"63820702",
        2152 => x"13050400",
        2153 => x"03248101",
        2154 => x"8320c101",
        2155 => x"83244101",
        2156 => x"03290101",
        2157 => x"8329c100",
        2158 => x"13010102",
        2159 => x"67800700",
        2160 => x"8320c101",
        2161 => x"03248101",
        2162 => x"83244101",
        2163 => x"03290101",
        2164 => x"8329c100",
        2165 => x"13010102",
        2166 => x"67800000",
        2167 => x"67800000",
        2168 => x"130101ff",
        2169 => x"23248100",
        2170 => x"23229100",
        2171 => x"93040500",
        2172 => x"13850500",
        2173 => x"93050600",
        2174 => x"13860600",
        2175 => x"23261100",
        2176 => x"23ac0186",
        2177 => x"ef10c057",
        2178 => x"9307f0ff",
        2179 => x"6318f500",
        2180 => x"83a78187",
        2181 => x"63840700",
        2182 => x"23a0f400",
        2183 => x"8320c100",
        2184 => x"03248100",
        2185 => x"83244100",
        2186 => x"13010101",
        2187 => x"67800000",
        2188 => x"130101ff",
        2189 => x"23248100",
        2190 => x"23229100",
        2191 => x"93040500",
        2192 => x"13850500",
        2193 => x"93050600",
        2194 => x"13860600",
        2195 => x"23261100",
        2196 => x"23ac0186",
        2197 => x"ef10c056",
        2198 => x"9307f0ff",
        2199 => x"6318f500",
        2200 => x"83a78187",
        2201 => x"63840700",
        2202 => x"23a0f400",
        2203 => x"8320c100",
        2204 => x"03248100",
        2205 => x"83244100",
        2206 => x"13010101",
        2207 => x"67800000",
        2208 => x"130101ff",
        2209 => x"23248100",
        2210 => x"23229100",
        2211 => x"93040500",
        2212 => x"13850500",
        2213 => x"93050600",
        2214 => x"13860600",
        2215 => x"23261100",
        2216 => x"23ac0186",
        2217 => x"ef10405c",
        2218 => x"9307f0ff",
        2219 => x"6318f500",
        2220 => x"83a78187",
        2221 => x"63840700",
        2222 => x"23a0f400",
        2223 => x"8320c100",
        2224 => x"03248100",
        2225 => x"83244100",
        2226 => x"13010101",
        2227 => x"67800000",
        2228 => x"03a50187",
        2229 => x"67800000",
        2230 => x"130101ff",
        2231 => x"23248100",
        2232 => x"23229100",
        2233 => x"37440000",
        2234 => x"b7440000",
        2235 => x"130444d8",
        2236 => x"938444d8",
        2237 => x"b3848440",
        2238 => x"23202101",
        2239 => x"23261100",
        2240 => x"93d42440",
        2241 => x"13090000",
        2242 => x"631e9902",
        2243 => x"37440000",
        2244 => x"b7440000",
        2245 => x"130444d8",
        2246 => x"938444d8",
        2247 => x"b3848440",
        2248 => x"93d42440",
        2249 => x"13090000",
        2250 => x"63189902",
        2251 => x"8320c100",
        2252 => x"03248100",
        2253 => x"83244100",
        2254 => x"03290100",
        2255 => x"13010101",
        2256 => x"67800000",
        2257 => x"83270400",
        2258 => x"13091900",
        2259 => x"13044400",
        2260 => x"e7800700",
        2261 => x"6ff05ffb",
        2262 => x"83270400",
        2263 => x"13091900",
        2264 => x"13044400",
        2265 => x"e7800700",
        2266 => x"6ff01ffc",
        2267 => x"13860500",
        2268 => x"93050500",
        2269 => x"03a50187",
        2270 => x"6f10801b",
        2271 => x"638a050e",
        2272 => x"83a7c5ff",
        2273 => x"130101fe",
        2274 => x"232c8100",
        2275 => x"232e1100",
        2276 => x"1384c5ff",
        2277 => x"63d40700",
        2278 => x"3304f400",
        2279 => x"2326a100",
        2280 => x"ef004031",
        2281 => x"83a70188",
        2282 => x"0325c100",
        2283 => x"639e0700",
        2284 => x"23220400",
        2285 => x"23a08188",
        2286 => x"03248101",
        2287 => x"8320c101",
        2288 => x"13010102",
        2289 => x"6f00402f",
        2290 => x"6374f402",
        2291 => x"03260400",
        2292 => x"b306c400",
        2293 => x"639ad700",
        2294 => x"83a60700",
        2295 => x"83a74700",
        2296 => x"b386c600",
        2297 => x"2320d400",
        2298 => x"2322f400",
        2299 => x"6ff09ffc",
        2300 => x"13870700",
        2301 => x"83a74700",
        2302 => x"63840700",
        2303 => x"e37af4fe",
        2304 => x"83260700",
        2305 => x"3306d700",
        2306 => x"63188602",
        2307 => x"03260400",
        2308 => x"b386c600",
        2309 => x"2320d700",
        2310 => x"3306d700",
        2311 => x"e39ec7f8",
        2312 => x"03a60700",
        2313 => x"83a74700",
        2314 => x"b306d600",
        2315 => x"2320d700",
        2316 => x"2322f700",
        2317 => x"6ff05ff8",
        2318 => x"6378c400",
        2319 => x"9307c000",
        2320 => x"2320f500",
        2321 => x"6ff05ff7",
        2322 => x"03260400",
        2323 => x"b306c400",
        2324 => x"639ad700",
        2325 => x"83a60700",
        2326 => x"83a74700",
        2327 => x"b386c600",
        2328 => x"2320d400",
        2329 => x"2322f400",
        2330 => x"23228700",
        2331 => x"6ff0dff4",
        2332 => x"67800000",
        2333 => x"130101ff",
        2334 => x"23248100",
        2335 => x"83a7c187",
        2336 => x"23229100",
        2337 => x"23202101",
        2338 => x"23261100",
        2339 => x"13090500",
        2340 => x"93840500",
        2341 => x"63980700",
        2342 => x"93050000",
        2343 => x"ef10000e",
        2344 => x"23aea186",
        2345 => x"93850400",
        2346 => x"13050900",
        2347 => x"ef10000d",
        2348 => x"9304f0ff",
        2349 => x"63129502",
        2350 => x"1304f0ff",
        2351 => x"8320c100",
        2352 => x"13050400",
        2353 => x"03248100",
        2354 => x"83244100",
        2355 => x"03290100",
        2356 => x"13010101",
        2357 => x"67800000",
        2358 => x"13043500",
        2359 => x"1374c4ff",
        2360 => x"e30e85fc",
        2361 => x"b305a440",
        2362 => x"13050900",
        2363 => x"ef100009",
        2364 => x"e31695fc",
        2365 => x"6ff05ffc",
        2366 => x"130101fe",
        2367 => x"232a9100",
        2368 => x"93843500",
        2369 => x"93f4c4ff",
        2370 => x"232e1100",
        2371 => x"232c8100",
        2372 => x"23282101",
        2373 => x"23263101",
        2374 => x"23244101",
        2375 => x"93848400",
        2376 => x"9307c000",
        2377 => x"63f4f400",
        2378 => x"93840700",
        2379 => x"63c40400",
        2380 => x"63f8b402",
        2381 => x"9307c000",
        2382 => x"2320f500",
        2383 => x"13050000",
        2384 => x"8320c101",
        2385 => x"03248101",
        2386 => x"83244101",
        2387 => x"03290101",
        2388 => x"8329c100",
        2389 => x"032a8100",
        2390 => x"13010102",
        2391 => x"67800000",
        2392 => x"13090500",
        2393 => x"ef000015",
        2394 => x"83a70188",
        2395 => x"13840700",
        2396 => x"63100408",
        2397 => x"93850400",
        2398 => x"13050900",
        2399 => x"eff09fef",
        2400 => x"9307f0ff",
        2401 => x"13040500",
        2402 => x"6312f512",
        2403 => x"03a40188",
        2404 => x"93070400",
        2405 => x"6392070e",
        2406 => x"63000410",
        2407 => x"032a0400",
        2408 => x"93050000",
        2409 => x"13050900",
        2410 => x"330a4401",
        2411 => x"ef00107d",
        2412 => x"6314aa0e",
        2413 => x"83270400",
        2414 => x"13050900",
        2415 => x"b384f440",
        2416 => x"93850400",
        2417 => x"eff01feb",
        2418 => x"9307f0ff",
        2419 => x"6306f50c",
        2420 => x"83270400",
        2421 => x"b3879700",
        2422 => x"2320f400",
        2423 => x"83a70188",
        2424 => x"03a74700",
        2425 => x"6310070a",
        2426 => x"23a00188",
        2427 => x"6f004003",
        2428 => x"83260400",
        2429 => x"b3869640",
        2430 => x"63ca0606",
        2431 => x"1307b000",
        2432 => x"637ad704",
        2433 => x"23209400",
        2434 => x"33079400",
        2435 => x"63908704",
        2436 => x"23a0e188",
        2437 => x"83274400",
        2438 => x"2320d700",
        2439 => x"2322f700",
        2440 => x"13050900",
        2441 => x"ef004009",
        2442 => x"1305b400",
        2443 => x"93074400",
        2444 => x"137585ff",
        2445 => x"3307f540",
        2446 => x"e304f5f0",
        2447 => x"3304e400",
        2448 => x"b387a740",
        2449 => x"2320f400",
        2450 => x"6ff09fef",
        2451 => x"23a2e700",
        2452 => x"6ff05ffc",
        2453 => x"03274400",
        2454 => x"63968700",
        2455 => x"23a0e188",
        2456 => x"6ff01ffc",
        2457 => x"23a2e700",
        2458 => x"6ff09ffb",
        2459 => x"93070400",
        2460 => x"03244400",
        2461 => x"6ff0dfef",
        2462 => x"13840700",
        2463 => x"83a74700",
        2464 => x"6ff05ff1",
        2465 => x"13870700",
        2466 => x"83a74700",
        2467 => x"e39c87fe",
        2468 => x"23220700",
        2469 => x"6ff0dff8",
        2470 => x"9307c000",
        2471 => x"2320f900",
        2472 => x"13050900",
        2473 => x"ef004001",
        2474 => x"6ff05fe9",
        2475 => x"23209500",
        2476 => x"6ff01ff7",
        2477 => x"67800000",
        2478 => x"67800000",
        2479 => x"130101fe",
        2480 => x"23282101",
        2481 => x"03a98500",
        2482 => x"232c8100",
        2483 => x"23263101",
        2484 => x"23206101",
        2485 => x"232e1100",
        2486 => x"232a9100",
        2487 => x"23244101",
        2488 => x"23225101",
        2489 => x"13840500",
        2490 => x"130b0600",
        2491 => x"93890600",
        2492 => x"63ec2613",
        2493 => x"8397c500",
        2494 => x"13070900",
        2495 => x"93f60748",
        2496 => x"638c0608",
        2497 => x"83244401",
        2498 => x"13073000",
        2499 => x"83a50501",
        2500 => x"b384e402",
        2501 => x"13072000",
        2502 => x"032a0400",
        2503 => x"930a0500",
        2504 => x"330aba40",
        2505 => x"b3c4e402",
        2506 => x"13871900",
        2507 => x"33074701",
        2508 => x"13860400",
        2509 => x"63f6e400",
        2510 => x"93040700",
        2511 => x"13060700",
        2512 => x"93f70740",
        2513 => x"6386070a",
        2514 => x"93050600",
        2515 => x"13850a00",
        2516 => x"eff09fda",
        2517 => x"13090500",
        2518 => x"630a050a",
        2519 => x"83250401",
        2520 => x"13060a00",
        2521 => x"efe09fc6",
        2522 => x"8357c400",
        2523 => x"93f7f7b7",
        2524 => x"93e70708",
        2525 => x"2316f400",
        2526 => x"23282401",
        2527 => x"232a9400",
        2528 => x"33094901",
        2529 => x"b3844441",
        2530 => x"23202401",
        2531 => x"23249400",
        2532 => x"13890900",
        2533 => x"13870900",
        2534 => x"93090700",
        2535 => x"03250400",
        2536 => x"13860900",
        2537 => x"93050b00",
        2538 => x"efe09fc4",
        2539 => x"83278400",
        2540 => x"13050000",
        2541 => x"b3872741",
        2542 => x"2324f400",
        2543 => x"83270400",
        2544 => x"b3873701",
        2545 => x"2320f400",
        2546 => x"8320c101",
        2547 => x"03248101",
        2548 => x"83244101",
        2549 => x"03290101",
        2550 => x"8329c100",
        2551 => x"032a8100",
        2552 => x"832a4100",
        2553 => x"032b0100",
        2554 => x"13010102",
        2555 => x"67800000",
        2556 => x"13850a00",
        2557 => x"ef00105d",
        2558 => x"13090500",
        2559 => x"e31e05f6",
        2560 => x"83250401",
        2561 => x"13850a00",
        2562 => x"eff05fb7",
        2563 => x"9307c000",
        2564 => x"23a0fa00",
        2565 => x"8357c400",
        2566 => x"1305f0ff",
        2567 => x"93e70704",
        2568 => x"2316f400",
        2569 => x"6ff05ffa",
        2570 => x"13890600",
        2571 => x"6ff01ff7",
        2572 => x"83278600",
        2573 => x"130101fd",
        2574 => x"232e3101",
        2575 => x"23261102",
        2576 => x"23248102",
        2577 => x"23229102",
        2578 => x"23202103",
        2579 => x"232c4101",
        2580 => x"232a5101",
        2581 => x"23286101",
        2582 => x"23267101",
        2583 => x"23248101",
        2584 => x"23229101",
        2585 => x"2320a101",
        2586 => x"93090600",
        2587 => x"63800710",
        2588 => x"032a0600",
        2589 => x"930c0500",
        2590 => x"13840500",
        2591 => x"930a3000",
        2592 => x"130b2000",
        2593 => x"83270a00",
        2594 => x"032c4a00",
        2595 => x"138d0700",
        2596 => x"630e0c10",
        2597 => x"03298400",
        2598 => x"93040900",
        2599 => x"636a2c15",
        2600 => x"8317c400",
        2601 => x"13f70748",
        2602 => x"63060708",
        2603 => x"83244401",
        2604 => x"83250401",
        2605 => x"832b0400",
        2606 => x"b3845403",
        2607 => x"b38bbb40",
        2608 => x"13871b00",
        2609 => x"33078701",
        2610 => x"b3c46403",
        2611 => x"13860400",
        2612 => x"63f6e400",
        2613 => x"93040700",
        2614 => x"13060700",
        2615 => x"93f70740",
        2616 => x"638a070c",
        2617 => x"93050600",
        2618 => x"13850c00",
        2619 => x"eff0dfc0",
        2620 => x"13090500",
        2621 => x"630e050c",
        2622 => x"83250401",
        2623 => x"13860b00",
        2624 => x"efe0dfac",
        2625 => x"8357c400",
        2626 => x"93f7f7b7",
        2627 => x"93e70708",
        2628 => x"2316f400",
        2629 => x"23282401",
        2630 => x"232a9400",
        2631 => x"33097901",
        2632 => x"b3847441",
        2633 => x"23202401",
        2634 => x"23249400",
        2635 => x"13090c00",
        2636 => x"93040c00",
        2637 => x"03250400",
        2638 => x"13860400",
        2639 => x"93050d00",
        2640 => x"efe01fab",
        2641 => x"83278400",
        2642 => x"b3872741",
        2643 => x"2324f400",
        2644 => x"83270400",
        2645 => x"b3879700",
        2646 => x"2320f400",
        2647 => x"83a78900",
        2648 => x"b3878741",
        2649 => x"23a4f900",
        2650 => x"63920704",
        2651 => x"13050000",
        2652 => x"8320c102",
        2653 => x"03248102",
        2654 => x"23a20900",
        2655 => x"83244102",
        2656 => x"03290102",
        2657 => x"8329c101",
        2658 => x"032a8101",
        2659 => x"832a4101",
        2660 => x"032b0101",
        2661 => x"832bc100",
        2662 => x"032c8100",
        2663 => x"832c4100",
        2664 => x"032d0100",
        2665 => x"13010103",
        2666 => x"67800000",
        2667 => x"130a8a00",
        2668 => x"6ff05fed",
        2669 => x"13850c00",
        2670 => x"ef00d040",
        2671 => x"13090500",
        2672 => x"e31a05f4",
        2673 => x"83250401",
        2674 => x"13850c00",
        2675 => x"eff01f9b",
        2676 => x"9307c000",
        2677 => x"23a0fc00",
        2678 => x"8357c400",
        2679 => x"1305f0ff",
        2680 => x"93e70704",
        2681 => x"2316f400",
        2682 => x"23a40900",
        2683 => x"6ff05ff8",
        2684 => x"13090c00",
        2685 => x"6ff0dff3",
        2686 => x"83d7c500",
        2687 => x"130101f5",
        2688 => x"2322910a",
        2689 => x"23248109",
        2690 => x"2326110a",
        2691 => x"2324810a",
        2692 => x"2320210b",
        2693 => x"232e3109",
        2694 => x"232c4109",
        2695 => x"232a5109",
        2696 => x"23286109",
        2697 => x"23267109",
        2698 => x"93f70708",
        2699 => x"130c0500",
        2700 => x"93840500",
        2701 => x"638a0706",
        2702 => x"83a70501",
        2703 => x"63960706",
        2704 => x"93050004",
        2705 => x"2326d100",
        2706 => x"2324c100",
        2707 => x"eff0dfaa",
        2708 => x"23a0a400",
        2709 => x"23a8a400",
        2710 => x"03268100",
        2711 => x"8326c100",
        2712 => x"63100504",
        2713 => x"9307c000",
        2714 => x"2320fc00",
        2715 => x"1305f0ff",
        2716 => x"8320c10a",
        2717 => x"0324810a",
        2718 => x"8324410a",
        2719 => x"0329010a",
        2720 => x"8329c109",
        2721 => x"032a8109",
        2722 => x"832a4109",
        2723 => x"032b0109",
        2724 => x"832bc108",
        2725 => x"032c8108",
        2726 => x"1301010b",
        2727 => x"67800000",
        2728 => x"93070004",
        2729 => x"23aaf400",
        2730 => x"93070002",
        2731 => x"a30cf102",
        2732 => x"b7490000",
        2733 => x"93070003",
        2734 => x"232a0102",
        2735 => x"230df102",
        2736 => x"232ed100",
        2737 => x"130af0ff",
        2738 => x"938909cf",
        2739 => x"130b1000",
        2740 => x"930aa000",
        2741 => x"13040600",
        2742 => x"83470400",
        2743 => x"b33bf000",
        2744 => x"9387b7fd",
        2745 => x"b337f000",
        2746 => x"b3fbfb00",
        2747 => x"63900b0c",
        2748 => x"b306c440",
        2749 => x"6304c402",
        2750 => x"93850400",
        2751 => x"13050c00",
        2752 => x"2324d100",
        2753 => x"eff09fbb",
        2754 => x"630c4523",
        2755 => x"83274103",
        2756 => x"83268100",
        2757 => x"b387d700",
        2758 => x"232af102",
        2759 => x"83470400",
        2760 => x"63800722",
        2761 => x"13041400",
        2762 => x"23200102",
        2763 => x"23260102",
        2764 => x"23224103",
        2765 => x"23240102",
        2766 => x"a3010106",
        2767 => x"232c0106",
        2768 => x"83450400",
        2769 => x"13065000",
        2770 => x"13850900",
        2771 => x"ef00101c",
        2772 => x"83270102",
        2773 => x"93061400",
        2774 => x"631e0504",
        2775 => x"13f70701",
        2776 => x"63060700",
        2777 => x"13070002",
        2778 => x"a301e106",
        2779 => x"13f78700",
        2780 => x"63060700",
        2781 => x"1307b002",
        2782 => x"a301e106",
        2783 => x"03460400",
        2784 => x"1307a002",
        2785 => x"6304e604",
        2786 => x"8327c102",
        2787 => x"93060000",
        2788 => x"13069000",
        2789 => x"03470400",
        2790 => x"130707fd",
        2791 => x"637ee608",
        2792 => x"63840604",
        2793 => x"2326f102",
        2794 => x"6f000004",
        2795 => x"13041400",
        2796 => x"6ff09ff2",
        2797 => x"33053541",
        2798 => x"3315ab00",
        2799 => x"3365f500",
        2800 => x"2320a102",
        2801 => x"13840600",
        2802 => x"6ff09ff7",
        2803 => x"0327c101",
        2804 => x"13064700",
        2805 => x"03270700",
        2806 => x"232ec100",
        2807 => x"63440704",
        2808 => x"2326e102",
        2809 => x"13840600",
        2810 => x"03470400",
        2811 => x"9307e002",
        2812 => x"631ef706",
        2813 => x"03471400",
        2814 => x"9307a002",
        2815 => x"6318f704",
        2816 => x"8327c101",
        2817 => x"13042400",
        2818 => x"13874700",
        2819 => x"83a70700",
        2820 => x"232ee100",
        2821 => x"63d40700",
        2822 => x"9307f0ff",
        2823 => x"2322f102",
        2824 => x"6f00c004",
        2825 => x"3307e040",
        2826 => x"93e72700",
        2827 => x"2326e102",
        2828 => x"2320f102",
        2829 => x"6ff01ffb",
        2830 => x"b3875703",
        2831 => x"13041400",
        2832 => x"93061000",
        2833 => x"b387e700",
        2834 => x"6ff0dff4",
        2835 => x"13041400",
        2836 => x"23220102",
        2837 => x"93070000",
        2838 => x"93069000",
        2839 => x"03470400",
        2840 => x"130707fd",
        2841 => x"63f8e608",
        2842 => x"e39a0bfa",
        2843 => x"83450400",
        2844 => x"b74b0000",
        2845 => x"13063000",
        2846 => x"13858bcf",
        2847 => x"ef001009",
        2848 => x"63020502",
        2849 => x"83270102",
        2850 => x"938b8bcf",
        2851 => x"33057541",
        2852 => x"13070004",
        2853 => x"3317a700",
        2854 => x"b3e7e700",
        2855 => x"13041400",
        2856 => x"2320f102",
        2857 => x"83450400",
        2858 => x"37450000",
        2859 => x"13066000",
        2860 => x"1305c5cf",
        2861 => x"230cb102",
        2862 => x"ef005005",
        2863 => x"630c0508",
        2864 => x"93070000",
        2865 => x"639a0704",
        2866 => x"03270102",
        2867 => x"8327c101",
        2868 => x"13770710",
        2869 => x"630a0702",
        2870 => x"93874700",
        2871 => x"232ef100",
        2872 => x"83274103",
        2873 => x"13061400",
        2874 => x"b3872701",
        2875 => x"232af102",
        2876 => x"6ff05fde",
        2877 => x"b3875703",
        2878 => x"13041400",
        2879 => x"930b1000",
        2880 => x"b387e700",
        2881 => x"6ff09ff5",
        2882 => x"93877700",
        2883 => x"93f787ff",
        2884 => x"93878700",
        2885 => x"6ff09ffc",
        2886 => x"b7260000",
        2887 => x"1307c101",
        2888 => x"9386c66b",
        2889 => x"13860400",
        2890 => x"93050102",
        2891 => x"13050c00",
        2892 => x"97000000",
        2893 => x"e7000000",
        2894 => x"13090500",
        2895 => x"e31245fb",
        2896 => x"83d7c400",
        2897 => x"93f70704",
        2898 => x"e39207d2",
        2899 => x"03254103",
        2900 => x"6ff01fd2",
        2901 => x"b7260000",
        2902 => x"1307c101",
        2903 => x"9386c66b",
        2904 => x"13860400",
        2905 => x"93050102",
        2906 => x"13050c00",
        2907 => x"ef00c01b",
        2908 => x"6ff09ffc",
        2909 => x"130101fd",
        2910 => x"232e3101",
        2911 => x"83a70501",
        2912 => x"93090700",
        2913 => x"03a78500",
        2914 => x"23248102",
        2915 => x"23202103",
        2916 => x"23286101",
        2917 => x"23267101",
        2918 => x"23261102",
        2919 => x"23229102",
        2920 => x"232c4101",
        2921 => x"232a5101",
        2922 => x"130b0500",
        2923 => x"13840500",
        2924 => x"13090600",
        2925 => x"938b0600",
        2926 => x"63d4e700",
        2927 => x"93070700",
        2928 => x"2320f900",
        2929 => x"03473404",
        2930 => x"63060700",
        2931 => x"93871700",
        2932 => x"2320f900",
        2933 => x"83270400",
        2934 => x"93f70702",
        2935 => x"63880700",
        2936 => x"83270900",
        2937 => x"93872700",
        2938 => x"2320f900",
        2939 => x"83240400",
        2940 => x"93f46400",
        2941 => x"639e0400",
        2942 => x"130a9401",
        2943 => x"930af0ff",
        2944 => x"8327c400",
        2945 => x"03270900",
        2946 => x"b387e740",
        2947 => x"63c4f408",
        2948 => x"83270400",
        2949 => x"83463404",
        2950 => x"93f70702",
        2951 => x"b336d000",
        2952 => x"6392070c",
        2953 => x"13063404",
        2954 => x"93850b00",
        2955 => x"13050b00",
        2956 => x"e7800900",
        2957 => x"9307f0ff",
        2958 => x"630af506",
        2959 => x"83270400",
        2960 => x"13074000",
        2961 => x"93040000",
        2962 => x"93f76700",
        2963 => x"639ee700",
        2964 => x"83270900",
        2965 => x"8324c400",
        2966 => x"b384f440",
        2967 => x"93c7f4ff",
        2968 => x"93d7f741",
        2969 => x"b3f4f400",
        2970 => x"83278400",
        2971 => x"03270401",
        2972 => x"6356f700",
        2973 => x"b387e740",
        2974 => x"b384f400",
        2975 => x"13090000",
        2976 => x"1304a401",
        2977 => x"130af0ff",
        2978 => x"63902409",
        2979 => x"13050000",
        2980 => x"6f000002",
        2981 => x"93061000",
        2982 => x"13060a00",
        2983 => x"93850b00",
        2984 => x"13050b00",
        2985 => x"e7800900",
        2986 => x"631a5503",
        2987 => x"1305f0ff",
        2988 => x"8320c102",
        2989 => x"03248102",
        2990 => x"83244102",
        2991 => x"03290102",
        2992 => x"8329c101",
        2993 => x"032a8101",
        2994 => x"832a4101",
        2995 => x"032b0101",
        2996 => x"832bc100",
        2997 => x"13010103",
        2998 => x"67800000",
        2999 => x"93841400",
        3000 => x"6ff01ff2",
        3001 => x"3307d400",
        3002 => x"13060003",
        3003 => x"a301c704",
        3004 => x"03475404",
        3005 => x"93871600",
        3006 => x"b307f400",
        3007 => x"93862600",
        3008 => x"a381e704",
        3009 => x"6ff01ff2",
        3010 => x"93061000",
        3011 => x"13060400",
        3012 => x"93850b00",
        3013 => x"13050b00",
        3014 => x"e7800900",
        3015 => x"e30845f9",
        3016 => x"13091900",
        3017 => x"6ff05ff6",
        3018 => x"130101fc",
        3019 => x"232c8102",
        3020 => x"232a9102",
        3021 => x"23244103",
        3022 => x"23225103",
        3023 => x"232e1102",
        3024 => x"23282103",
        3025 => x"23263103",
        3026 => x"83c78501",
        3027 => x"93840600",
        3028 => x"93068007",
        3029 => x"130a0500",
        3030 => x"13840500",
        3031 => x"930a0600",
        3032 => x"63eef600",
        3033 => x"93062006",
        3034 => x"13863504",
        3035 => x"63ecf600",
        3036 => x"63820728",
        3037 => x"93068005",
        3038 => x"638ed720",
        3039 => x"13092404",
        3040 => x"6f000004",
        3041 => x"9386d7f9",
        3042 => x"93f6f60f",
        3043 => x"93055001",
        3044 => x"e3e6d5fe",
        3045 => x"b7450000",
        3046 => x"93962600",
        3047 => x"9385c5d2",
        3048 => x"b386b600",
        3049 => x"83a60600",
        3050 => x"67800600",
        3051 => x"83270700",
        3052 => x"13092404",
        3053 => x"93864700",
        3054 => x"83a70700",
        3055 => x"2320d700",
        3056 => x"2301f404",
        3057 => x"93071000",
        3058 => x"6f008026",
        3059 => x"83270400",
        3060 => x"03250700",
        3061 => x"93f60708",
        3062 => x"93054500",
        3063 => x"63860602",
        3064 => x"83270500",
        3065 => x"2320b700",
        3066 => x"b7460000",
        3067 => x"63d80700",
        3068 => x"1307d002",
        3069 => x"b307f040",
        3070 => x"a301e404",
        3071 => x"938646d0",
        3072 => x"1307a000",
        3073 => x"6f008006",
        3074 => x"93f60704",
        3075 => x"83270500",
        3076 => x"2320b700",
        3077 => x"e38a06fc",
        3078 => x"93970701",
        3079 => x"93d70741",
        3080 => x"6ff09ffc",
        3081 => x"83250400",
        3082 => x"83260700",
        3083 => x"13f50508",
        3084 => x"83a70600",
        3085 => x"93864600",
        3086 => x"631a0500",
        3087 => x"93f50504",
        3088 => x"63860500",
        3089 => x"93970701",
        3090 => x"93d70701",
        3091 => x"2320d700",
        3092 => x"83458401",
        3093 => x"b7460000",
        3094 => x"1307f006",
        3095 => x"938646d0",
        3096 => x"6398e514",
        3097 => x"13078000",
        3098 => x"a3010404",
        3099 => x"83254400",
        3100 => x"2324b400",
        3101 => x"63ce0500",
        3102 => x"03250400",
        3103 => x"b3e5b700",
        3104 => x"13090600",
        3105 => x"1375b5ff",
        3106 => x"2320a400",
        3107 => x"63840502",
        3108 => x"13090600",
        3109 => x"b3f5e702",
        3110 => x"1309f9ff",
        3111 => x"b385b600",
        3112 => x"83c50500",
        3113 => x"2300b900",
        3114 => x"93850700",
        3115 => x"b3d7e702",
        3116 => x"e3f2e5fe",
        3117 => x"93078000",
        3118 => x"6314f702",
        3119 => x"83270400",
        3120 => x"93f71700",
        3121 => x"638e0700",
        3122 => x"03274400",
        3123 => x"83270401",
        3124 => x"63c8e700",
        3125 => x"93070003",
        3126 => x"a30ff9fe",
        3127 => x"1309f9ff",
        3128 => x"33062641",
        3129 => x"2328c400",
        3130 => x"13870400",
        3131 => x"93860a00",
        3132 => x"1306c101",
        3133 => x"93050400",
        3134 => x"13050a00",
        3135 => x"eff09fc7",
        3136 => x"9309f0ff",
        3137 => x"631c3513",
        3138 => x"1305f0ff",
        3139 => x"8320c103",
        3140 => x"03248103",
        3141 => x"83244103",
        3142 => x"03290103",
        3143 => x"8329c102",
        3144 => x"032a8102",
        3145 => x"832a4102",
        3146 => x"13010104",
        3147 => x"67800000",
        3148 => x"83270400",
        3149 => x"93e70702",
        3150 => x"2320f400",
        3151 => x"b7460000",
        3152 => x"93078007",
        3153 => x"938686d1",
        3154 => x"a302f404",
        3155 => x"83250400",
        3156 => x"03250700",
        3157 => x"13f80508",
        3158 => x"83270500",
        3159 => x"13054500",
        3160 => x"631a0800",
        3161 => x"13f80504",
        3162 => x"63060800",
        3163 => x"93970701",
        3164 => x"93d70701",
        3165 => x"2320a700",
        3166 => x"13f71500",
        3167 => x"63060700",
        3168 => x"93e50502",
        3169 => x"2320b400",
        3170 => x"638c0700",
        3171 => x"13070001",
        3172 => x"6ff09fed",
        3173 => x"b7460000",
        3174 => x"938646d0",
        3175 => x"6ff0dffa",
        3176 => x"03270400",
        3177 => x"1377f7fd",
        3178 => x"2320e400",
        3179 => x"6ff01ffe",
        3180 => x"1307a000",
        3181 => x"6ff05feb",
        3182 => x"83260400",
        3183 => x"83270700",
        3184 => x"83254401",
        3185 => x"13f80608",
        3186 => x"13854700",
        3187 => x"630a0800",
        3188 => x"2320a700",
        3189 => x"83a70700",
        3190 => x"23a0b700",
        3191 => x"6f008001",
        3192 => x"2320a700",
        3193 => x"93f60604",
        3194 => x"83a70700",
        3195 => x"e38606fe",
        3196 => x"2390b700",
        3197 => x"23280400",
        3198 => x"13090600",
        3199 => x"6ff0dfee",
        3200 => x"83270700",
        3201 => x"03264400",
        3202 => x"93050000",
        3203 => x"93864700",
        3204 => x"2320d700",
        3205 => x"03a90700",
        3206 => x"13050900",
        3207 => x"ef00002f",
        3208 => x"63060500",
        3209 => x"33052541",
        3210 => x"2322a400",
        3211 => x"83274400",
        3212 => x"2328f400",
        3213 => x"a3010404",
        3214 => x"6ff01feb",
        3215 => x"83260401",
        3216 => x"13060900",
        3217 => x"93850a00",
        3218 => x"13050a00",
        3219 => x"e7800400",
        3220 => x"e30c35eb",
        3221 => x"83270400",
        3222 => x"93f72700",
        3223 => x"63960704",
        3224 => x"8327c101",
        3225 => x"0325c400",
        3226 => x"e352f5ea",
        3227 => x"13850700",
        3228 => x"6ff0dfe9",
        3229 => x"93061000",
        3230 => x"93850a00",
        3231 => x"13050a00",
        3232 => x"2326c100",
        3233 => x"e7800400",
        3234 => x"e30035e9",
        3235 => x"0326c100",
        3236 => x"13091900",
        3237 => x"8327c400",
        3238 => x"0327c101",
        3239 => x"b387e740",
        3240 => x"e34af9fc",
        3241 => x"6ff0dffb",
        3242 => x"13090000",
        3243 => x"13069401",
        3244 => x"6ff05ffe",
        3245 => x"8397c500",
        3246 => x"130101fe",
        3247 => x"232c8100",
        3248 => x"232a9100",
        3249 => x"232e1100",
        3250 => x"23282101",
        3251 => x"13f78700",
        3252 => x"93040500",
        3253 => x"13840500",
        3254 => x"63120712",
        3255 => x"03a74500",
        3256 => x"6346e000",
        3257 => x"03a70504",
        3258 => x"6356e010",
        3259 => x"0327c402",
        3260 => x"63020710",
        3261 => x"03a90400",
        3262 => x"93963701",
        3263 => x"23a00400",
        3264 => x"63dc060a",
        3265 => x"03264405",
        3266 => x"8357c400",
        3267 => x"93f74700",
        3268 => x"638e0700",
        3269 => x"83274400",
        3270 => x"3306f640",
        3271 => x"83274403",
        3272 => x"63860700",
        3273 => x"83270404",
        3274 => x"3306f640",
        3275 => x"8327c402",
        3276 => x"83250402",
        3277 => x"93060000",
        3278 => x"13850400",
        3279 => x"e7800700",
        3280 => x"1307f0ff",
        3281 => x"8317c400",
        3282 => x"6312e502",
        3283 => x"83a60400",
        3284 => x"1307d001",
        3285 => x"636cd70e",
        3286 => x"37074020",
        3287 => x"13071700",
        3288 => x"3357d700",
        3289 => x"13771700",
        3290 => x"6302070e",
        3291 => x"03270401",
        3292 => x"23220400",
        3293 => x"2320e400",
        3294 => x"13973701",
        3295 => x"635c0700",
        3296 => x"9307f0ff",
        3297 => x"6316f500",
        3298 => x"83a70400",
        3299 => x"63940700",
        3300 => x"232aa404",
        3301 => x"83254403",
        3302 => x"23a02401",
        3303 => x"638c0504",
        3304 => x"93074404",
        3305 => x"6386f500",
        3306 => x"13850400",
        3307 => x"efe01ffd",
        3308 => x"232a0402",
        3309 => x"6f000004",
        3310 => x"83250402",
        3311 => x"13060000",
        3312 => x"93061000",
        3313 => x"13850400",
        3314 => x"e7000700",
        3315 => x"9307f0ff",
        3316 => x"13060500",
        3317 => x"e31af5f2",
        3318 => x"83a70400",
        3319 => x"e38607f2",
        3320 => x"138737fe",
        3321 => x"63060700",
        3322 => x"9387a7fe",
        3323 => x"639e0704",
        3324 => x"23a02401",
        3325 => x"13050000",
        3326 => x"6f000006",
        3327 => x"03a60501",
        3328 => x"e30a06fe",
        3329 => x"83a60500",
        3330 => x"93f73700",
        3331 => x"23a0c500",
        3332 => x"3389c640",
        3333 => x"13070000",
        3334 => x"63940700",
        3335 => x"03a74501",
        3336 => x"2324e400",
        3337 => x"e35820fd",
        3338 => x"83278402",
        3339 => x"83250402",
        3340 => x"93060900",
        3341 => x"13850400",
        3342 => x"2326c100",
        3343 => x"e7800700",
        3344 => x"0326c100",
        3345 => x"6346a002",
        3346 => x"8357c400",
        3347 => x"93e70704",
        3348 => x"2316f400",
        3349 => x"1305f0ff",
        3350 => x"8320c101",
        3351 => x"03248101",
        3352 => x"83244101",
        3353 => x"03290101",
        3354 => x"13010102",
        3355 => x"67800000",
        3356 => x"3306a600",
        3357 => x"3309a940",
        3358 => x"6ff0dffa",
        3359 => x"83a70501",
        3360 => x"638e0704",
        3361 => x"130101fe",
        3362 => x"232c8100",
        3363 => x"232e1100",
        3364 => x"13040500",
        3365 => x"630c0500",
        3366 => x"83270502",
        3367 => x"63980700",
        3368 => x"2326b100",
        3369 => x"efe09f86",
        3370 => x"8325c100",
        3371 => x"8397c500",
        3372 => x"638c0700",
        3373 => x"13050400",
        3374 => x"03248101",
        3375 => x"8320c101",
        3376 => x"13010102",
        3377 => x"6ff01fdf",
        3378 => x"8320c101",
        3379 => x"03248101",
        3380 => x"13050000",
        3381 => x"13010102",
        3382 => x"67800000",
        3383 => x"13050000",
        3384 => x"67800000",
        3385 => x"93050500",
        3386 => x"631e0500",
        3387 => x"b7350000",
        3388 => x"37050020",
        3389 => x"13868181",
        3390 => x"9385c547",
        3391 => x"13054502",
        3392 => x"6fe01f86",
        3393 => x"03a50187",
        3394 => x"6ff05ff7",
        3395 => x"93f5f50f",
        3396 => x"3306c500",
        3397 => x"6316c500",
        3398 => x"13050000",
        3399 => x"67800000",
        3400 => x"83470500",
        3401 => x"e38cb7fe",
        3402 => x"13051500",
        3403 => x"6ff09ffe",
        3404 => x"130101ff",
        3405 => x"23248100",
        3406 => x"23229100",
        3407 => x"93040500",
        3408 => x"13850500",
        3409 => x"93050600",
        3410 => x"23261100",
        3411 => x"23ac0186",
        3412 => x"ef00c01b",
        3413 => x"9307f0ff",
        3414 => x"6318f500",
        3415 => x"83a78187",
        3416 => x"63840700",
        3417 => x"23a0f400",
        3418 => x"8320c100",
        3419 => x"03248100",
        3420 => x"83244100",
        3421 => x"13010101",
        3422 => x"67800000",
        3423 => x"130101ff",
        3424 => x"23248100",
        3425 => x"23229100",
        3426 => x"93040500",
        3427 => x"13850500",
        3428 => x"23261100",
        3429 => x"23ac0186",
        3430 => x"ef008026",
        3431 => x"9307f0ff",
        3432 => x"6318f500",
        3433 => x"83a78187",
        3434 => x"63840700",
        3435 => x"23a0f400",
        3436 => x"8320c100",
        3437 => x"03248100",
        3438 => x"83244100",
        3439 => x"13010101",
        3440 => x"67800000",
        3441 => x"63960500",
        3442 => x"93050600",
        3443 => x"6fe0dff2",
        3444 => x"130101fe",
        3445 => x"232c8100",
        3446 => x"23244101",
        3447 => x"232e1100",
        3448 => x"232a9100",
        3449 => x"23282101",
        3450 => x"23263101",
        3451 => x"13040600",
        3452 => x"130a0500",
        3453 => x"63180602",
        3454 => x"efe05fd8",
        3455 => x"93040000",
        3456 => x"8320c101",
        3457 => x"03248101",
        3458 => x"03290101",
        3459 => x"8329c100",
        3460 => x"032a8100",
        3461 => x"13850400",
        3462 => x"83244101",
        3463 => x"13010102",
        3464 => x"67800000",
        3465 => x"93840500",
        3466 => x"ef008005",
        3467 => x"13090500",
        3468 => x"63668500",
        3469 => x"93571500",
        3470 => x"e3e487fc",
        3471 => x"93050400",
        3472 => x"13050a00",
        3473 => x"efe05feb",
        3474 => x"93090500",
        3475 => x"63160500",
        3476 => x"93840900",
        3477 => x"6ff0dffa",
        3478 => x"13060400",
        3479 => x"63748900",
        3480 => x"13060900",
        3481 => x"93850400",
        3482 => x"13850900",
        3483 => x"efd01fd6",
        3484 => x"93850400",
        3485 => x"13050a00",
        3486 => x"efe05fd0",
        3487 => x"6ff05ffd",
        3488 => x"83a7c5ff",
        3489 => x"1385c7ff",
        3490 => x"63d80700",
        3491 => x"b385a500",
        3492 => x"83a70500",
        3493 => x"3305f500",
        3494 => x"67800000",
        3495 => x"130101ff",
        3496 => x"23261100",
        3497 => x"23248100",
        3498 => x"93089003",
        3499 => x"73000000",
        3500 => x"13040500",
        3501 => x"635a0500",
        3502 => x"33048040",
        3503 => x"efe05fc1",
        3504 => x"23208500",
        3505 => x"1304f0ff",
        3506 => x"8320c100",
        3507 => x"13050400",
        3508 => x"03248100",
        3509 => x"13010101",
        3510 => x"67800000",
        3511 => x"9308d005",
        3512 => x"73000000",
        3513 => x"63520502",
        3514 => x"130101ff",
        3515 => x"23248100",
        3516 => x"13040500",
        3517 => x"23261100",
        3518 => x"33048040",
        3519 => x"efe05fbd",
        3520 => x"23208500",
        3521 => x"6f000000",
        3522 => x"6f000000",
        3523 => x"130101fe",
        3524 => x"232a9100",
        3525 => x"232e1100",
        3526 => x"93040500",
        3527 => x"232c8100",
        3528 => x"93083019",
        3529 => x"13050000",
        3530 => x"93050100",
        3531 => x"73000000",
        3532 => x"13040500",
        3533 => x"635a0500",
        3534 => x"33048040",
        3535 => x"efe05fb9",
        3536 => x"23208500",
        3537 => x"1304f0ff",
        3538 => x"83274100",
        3539 => x"03270100",
        3540 => x"8320c101",
        3541 => x"23a2f400",
        3542 => x"83278100",
        3543 => x"23a0e400",
        3544 => x"1307803e",
        3545 => x"b3c7e702",
        3546 => x"13050400",
        3547 => x"03248101",
        3548 => x"23a4f400",
        3549 => x"83244101",
        3550 => x"13010102",
        3551 => x"67800000",
        3552 => x"130101ff",
        3553 => x"23261100",
        3554 => x"23248100",
        3555 => x"9308e003",
        3556 => x"73000000",
        3557 => x"13040500",
        3558 => x"635a0500",
        3559 => x"33048040",
        3560 => x"efe01fb3",
        3561 => x"23208500",
        3562 => x"1304f0ff",
        3563 => x"8320c100",
        3564 => x"13050400",
        3565 => x"03248100",
        3566 => x"13010101",
        3567 => x"67800000",
        3568 => x"130101ff",
        3569 => x"23261100",
        3570 => x"23248100",
        3571 => x"9308f003",
        3572 => x"73000000",
        3573 => x"13040500",
        3574 => x"635a0500",
        3575 => x"33048040",
        3576 => x"efe01faf",
        3577 => x"23208500",
        3578 => x"1304f0ff",
        3579 => x"8320c100",
        3580 => x"13050400",
        3581 => x"03248100",
        3582 => x"13010101",
        3583 => x"67800000",
        3584 => x"93060500",
        3585 => x"03a54188",
        3586 => x"130101ff",
        3587 => x"23261100",
        3588 => x"631a0502",
        3589 => x"9308600d",
        3590 => x"73000000",
        3591 => x"9307f0ff",
        3592 => x"6310f502",
        3593 => x"efe0dfaa",
        3594 => x"9307c000",
        3595 => x"2320f500",
        3596 => x"1305f0ff",
        3597 => x"8320c100",
        3598 => x"13010101",
        3599 => x"67800000",
        3600 => x"23a2a188",
        3601 => x"9308600d",
        3602 => x"3385a600",
        3603 => x"73000000",
        3604 => x"83a74188",
        3605 => x"b386f600",
        3606 => x"e316d5fc",
        3607 => x"23a2a188",
        3608 => x"13850700",
        3609 => x"6ff01ffd",
        3610 => x"130101ff",
        3611 => x"23261100",
        3612 => x"23248100",
        3613 => x"93080004",
        3614 => x"73000000",
        3615 => x"13040500",
        3616 => x"635a0500",
        3617 => x"33048040",
        3618 => x"efe09fa4",
        3619 => x"23208500",
        3620 => x"1304f0ff",
        3621 => x"8320c100",
        3622 => x"13050400",
        3623 => x"03248100",
        3624 => x"13010101",
        3625 => x"67800000",
        3626 => x"10000000",
        3627 => x"00000000",
        3628 => x"037a5200",
        3629 => x"017c0101",
        3630 => x"1b0c0200",
        3631 => x"10000000",
        3632 => x"18000000",
        3633 => x"d8ceffff",
        3634 => x"0c040000",
        3635 => x"00000000",
        3636 => x"10000000",
        3637 => x"00000000",
        3638 => x"037a5200",
        3639 => x"017c0101",
        3640 => x"1b0c0200",
        3641 => x"10000000",
        3642 => x"18000000",
        3643 => x"bcd2ffff",
        3644 => x"ec030000",
        3645 => x"00000000",
        3646 => x"10000000",
        3647 => x"00000000",
        3648 => x"037a5200",
        3649 => x"017c0101",
        3650 => x"1b0c0200",
        3651 => x"10000000",
        3652 => x"18000000",
        3653 => x"80d6ffff",
        3654 => x"1c040000",
        3655 => x"00000000",
        3656 => x"30313233",
        3657 => x"34353637",
        3658 => x"38396162",
        3659 => x"63646566",
        3660 => x"00000000",
        3661 => x"a0040000",
        3662 => x"a4040000",
        3663 => x"a4040000",
        3664 => x"a4040000",
        3665 => x"14050000",
        3666 => x"a4040000",
        3667 => x"a4040000",
        3668 => x"a4040000",
        3669 => x"a4040000",
        3670 => x"a4040000",
        3671 => x"a4040000",
        3672 => x"a4040000",
        3673 => x"a4040000",
        3674 => x"a4040000",
        3675 => x"a4040000",
        3676 => x"1c050000",
        3677 => x"a4040000",
        3678 => x"34050000",
        3679 => x"3c050000",
        3680 => x"a4040000",
        3681 => x"44050000",
        3682 => x"4c050000",
        3683 => x"a4040000",
        3684 => x"24050000",
        3685 => x"2c050000",
        3686 => x"a0050000",
        3687 => x"80050000",
        3688 => x"80050000",
        3689 => x"80050000",
        3690 => x"80050000",
        3691 => x"a4040000",
        3692 => x"24060000",
        3693 => x"f0050000",
        3694 => x"80050000",
        3695 => x"80050000",
        3696 => x"80050000",
        3697 => x"80050000",
        3698 => x"80050000",
        3699 => x"80050000",
        3700 => x"80050000",
        3701 => x"80050000",
        3702 => x"80050000",
        3703 => x"80050000",
        3704 => x"80050000",
        3705 => x"80050000",
        3706 => x"80050000",
        3707 => x"80050000",
        3708 => x"94050000",
        3709 => x"94050000",
        3710 => x"80050000",
        3711 => x"80050000",
        3712 => x"80050000",
        3713 => x"80050000",
        3714 => x"80050000",
        3715 => x"80050000",
        3716 => x"80050000",
        3717 => x"80050000",
        3718 => x"80050000",
        3719 => x"80050000",
        3720 => x"80050000",
        3721 => x"80050000",
        3722 => x"a4040000",
        3723 => x"a0050000",
        3724 => x"b4050000",
        3725 => x"dc050000",
        3726 => x"80050000",
        3727 => x"80050000",
        3728 => x"80050000",
        3729 => x"80050000",
        3730 => x"80050000",
        3731 => x"80050000",
        3732 => x"c8050000",
        3733 => x"80050000",
        3734 => x"80050000",
        3735 => x"80050000",
        3736 => x"80050000",
        3737 => x"94050000",
        3738 => x"94050000",
        3739 => x"00010202",
        3740 => x"03030303",
        3741 => x"04040404",
        3742 => x"04040404",
        3743 => x"05050505",
        3744 => x"05050505",
        3745 => x"05050505",
        3746 => x"05050505",
        3747 => x"06060606",
        3748 => x"06060606",
        3749 => x"06060606",
        3750 => x"06060606",
        3751 => x"06060606",
        3752 => x"06060606",
        3753 => x"06060606",
        3754 => x"06060606",
        3755 => x"07070707",
        3756 => x"07070707",
        3757 => x"07070707",
        3758 => x"07070707",
        3759 => x"07070707",
        3760 => x"07070707",
        3761 => x"07070707",
        3762 => x"07070707",
        3763 => x"07070707",
        3764 => x"07070707",
        3765 => x"07070707",
        3766 => x"07070707",
        3767 => x"07070707",
        3768 => x"07070707",
        3769 => x"07070707",
        3770 => x"07070707",
        3771 => x"08080808",
        3772 => x"08080808",
        3773 => x"08080808",
        3774 => x"08080808",
        3775 => x"08080808",
        3776 => x"08080808",
        3777 => x"08080808",
        3778 => x"08080808",
        3779 => x"08080808",
        3780 => x"08080808",
        3781 => x"08080808",
        3782 => x"08080808",
        3783 => x"08080808",
        3784 => x"08080808",
        3785 => x"08080808",
        3786 => x"08080808",
        3787 => x"08080808",
        3788 => x"08080808",
        3789 => x"08080808",
        3790 => x"08080808",
        3791 => x"08080808",
        3792 => x"08080808",
        3793 => x"08080808",
        3794 => x"08080808",
        3795 => x"08080808",
        3796 => x"08080808",
        3797 => x"08080808",
        3798 => x"08080808",
        3799 => x"08080808",
        3800 => x"08080808",
        3801 => x"08080808",
        3802 => x"08080808",
        3803 => x"0d0a4542",
        3804 => x"5245414b",
        3805 => x"21206d65",
        3806 => x"7063203d",
        3807 => x"20000000",
        3808 => x"20696e73",
        3809 => x"6e203d20",
        3810 => x"00000000",
        3811 => x"0d0a0000",
        3812 => x"0d0a436c",
        3813 => x"6f636b20",
        3814 => x"66726571",
        3815 => x"75656e63",
        3816 => x"793a2000",
        3817 => x"0d0a4861",
        3818 => x"72647761",
        3819 => x"72652076",
        3820 => x"65727369",
        3821 => x"6f6e3a20",
        3822 => x"00000000",
        3823 => x"0d0a0a44",
        3824 => x"6973706c",
        3825 => x"6179696e",
        3826 => x"67207468",
        3827 => x"65207469",
        3828 => x"6d652070",
        3829 => x"61737365",
        3830 => x"64207369",
        3831 => x"6e636520",
        3832 => x"72657365",
        3833 => x"740d0a0a",
        3834 => x"00000000",
        3835 => x"4f6e2d63",
        3836 => x"68697020",
        3837 => x"64656275",
        3838 => x"67676572",
        3839 => x"20666f75",
        3840 => x"6e642c20",
        3841 => x"736b6970",
        3842 => x"70696e67",
        3843 => x"20454252",
        3844 => x"45414b20",
        3845 => x"696e7374",
        3846 => x"72756374",
        3847 => x"696f6e0d",
        3848 => x"0a0d0a00",
        3849 => x"2530356c",
        3850 => x"643a2530",
        3851 => x"366c6420",
        3852 => x"20202530",
        3853 => x"326c643a",
        3854 => x"2530326c",
        3855 => x"643a2530",
        3856 => x"326c640d",
        3857 => x"00000000",
        3858 => x"696e7465",
        3859 => x"72727570",
        3860 => x"745f6469",
        3861 => x"72656374",
        3862 => x"00000000",
        3863 => x"54485541",
        3864 => x"53205249",
        3865 => x"53432d56",
        3866 => x"20525633",
        3867 => x"32494d20",
        3868 => x"62617265",
        3869 => x"206d6574",
        3870 => x"616c2070",
        3871 => x"726f6365",
        3872 => x"73736f72",
        3873 => x"00000000",
        3874 => x"54686520",
        3875 => x"48616775",
        3876 => x"6520556e",
        3877 => x"69766572",
        3878 => x"73697479",
        3879 => x"206f6620",
        3880 => x"4170706c",
        3881 => x"69656420",
        3882 => x"53636965",
        3883 => x"6e636573",
        3884 => x"00000000",
        3885 => x"44657061",
        3886 => x"72746d65",
        3887 => x"6e74206f",
        3888 => x"6620456c",
        3889 => x"65637472",
        3890 => x"6963616c",
        3891 => x"20456e67",
        3892 => x"696e6565",
        3893 => x"72696e67",
        3894 => x"00000000",
        3895 => x"4a2e452e",
        3896 => x"4a2e206f",
        3897 => x"70206465",
        3898 => x"6e204272",
        3899 => x"6f757700",
        3900 => x"232d302b",
        3901 => x"20000000",
        3902 => x"686c4c00",
        3903 => x"65666745",
        3904 => x"46470000",
        3905 => x"30313233",
        3906 => x"34353637",
        3907 => x"38394142",
        3908 => x"43444546",
        3909 => x"00000000",
        3910 => x"30313233",
        3911 => x"34353637",
        3912 => x"38396162",
        3913 => x"63646566",
        3914 => x"00000000",
        3915 => x"ac2f0000",
        3916 => x"cc2f0000",
        3917 => x"7c2f0000",
        3918 => x"7c2f0000",
        3919 => x"7c2f0000",
        3920 => x"7c2f0000",
        3921 => x"cc2f0000",
        3922 => x"7c2f0000",
        3923 => x"7c2f0000",
        3924 => x"7c2f0000",
        3925 => x"7c2f0000",
        3926 => x"b8310000",
        3927 => x"24300000",
        3928 => x"30310000",
        3929 => x"7c2f0000",
        3930 => x"7c2f0000",
        3931 => x"00320000",
        3932 => x"7c2f0000",
        3933 => x"24300000",
        3934 => x"7c2f0000",
        3935 => x"7c2f0000",
        3936 => x"3c310000",
        3937 => x"483c0000",
        3938 => x"5c3c0000",
        3939 => x"883c0000",
        3940 => x"b43c0000",
        3941 => x"dc3c0000",
        3942 => x"00000000",
        3943 => x"00000000",
        3944 => x"03000000",
        3945 => x"88000020",
        3946 => x"00000000",
        3947 => x"88000020",
        3948 => x"f0000020",
        3949 => x"58010020",
        3950 => x"00000000",
        3951 => x"00000000",
        3952 => x"00000000",
        3953 => x"00000000",
        3954 => x"00000000",
        3955 => x"00000000",
        3956 => x"00000000",
        3957 => x"00000000",
        3958 => x"00000000",
        3959 => x"00000000",
        3960 => x"00000000",
        3961 => x"00000000",
        3962 => x"00000000",
        3963 => x"00000000",
        3964 => x"00000000",
        3965 => x"24000020"
            );
end package rom_image;
