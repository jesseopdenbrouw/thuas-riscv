-- srec2vhdl table generator
-- for input file 'bootloader.srec'
-- date: Sat Sep 13 23:13:30 2025


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package bootrom_image is
    constant bootrom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382826e",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"37060020",
           9 => x"13050500",
          10 => x"13060600",
          11 => x"637ac500",
          12 => x"b7150010",
          13 => x"3306a640",
          14 => x"938545f5",
          15 => x"ef00c06c",
          16 => x"37050020",
          17 => x"37060020",
          18 => x"13050500",
          19 => x"13060600",
          20 => x"6378c500",
          21 => x"3306a640",
          22 => x"93050000",
          23 => x"ef000069",
          24 => x"37c50100",
          25 => x"93051000",
          26 => x"13050520",
          27 => x"ef009007",
          28 => x"ef001039",
          29 => x"37150010",
          30 => x"130545de",
          31 => x"ef00900b",
          32 => x"732530f1",
          33 => x"93058000",
          34 => x"ef009030",
          35 => x"37150010",
          36 => x"130545e1",
          37 => x"ef00100a",
          38 => x"732510fc",
          39 => x"371a0010",
          40 => x"ef009024",
          41 => x"1305cad5",
          42 => x"ef00d008",
          43 => x"b70900f0",
          44 => x"9307f03f",
          45 => x"3709a000",
          46 => x"23a2f900",
          47 => x"13091900",
          48 => x"93041000",
          49 => x"6f008001",
          50 => x"ef00d000",
          51 => x"13040500",
          52 => x"93841400",
          53 => x"631a0502",
          54 => x"638e242b",
          55 => x"9397c400",
          56 => x"e39407fe",
          57 => x"1305a002",
          58 => x"ef00d002",
          59 => x"83a74900",
          60 => x"93841400",
          61 => x"93d71700",
          62 => x"23a2f900",
          63 => x"ef00807d",
          64 => x"13040500",
          65 => x"e30a05fc",
          66 => x"b70700f0",
          67 => x"23a20700",
          68 => x"ef00c061",
          69 => x"9377f50f",
          70 => x"13071002",
          71 => x"638ee744",
          72 => x"13074002",
          73 => x"6384e728",
          74 => x"232c0100",
          75 => x"97020000",
          76 => x"9382824e",
          77 => x"73905230",
          78 => x"1305cad5",
          79 => x"ef00807f",
          80 => x"b71a0010",
          81 => x"1387cae2",
          82 => x"2326e100",
          83 => x"b7770000",
          84 => x"37770000",
          85 => x"b7190010",
          86 => x"13072777",
          87 => x"93877777",
          88 => x"130acad5",
          89 => x"938999c5",
          90 => x"2328e100",
          91 => x"232af100",
          92 => x"13040000",
          93 => x"130b8006",
          94 => x"130d2007",
          95 => x"0325c100",
          96 => x"ef00407b",
          97 => x"13054102",
          98 => x"93059002",
          99 => x"ef00005c",
         100 => x"83574102",
         101 => x"93040500",
         102 => x"63806713",
         103 => x"6388a713",
         104 => x"03270101",
         105 => x"638ae714",
         106 => x"83574102",
         107 => x"03274101",
         108 => x"6384e71a",
         109 => x"03574102",
         110 => x"b7770000",
         111 => x"93874776",
         112 => x"630af702",
         113 => x"93071000",
         114 => x"03474102",
         115 => x"63800704",
         116 => x"9307e006",
         117 => x"6308f704",
         118 => x"e38204fa",
         119 => x"b7170010",
         120 => x"138507f5",
         121 => x"ef000075",
         122 => x"13050a00",
         123 => x"ef008074",
         124 => x"6ff0dff8",
         125 => x"03476102",
         126 => x"93070002",
         127 => x"e314f7fc",
         128 => x"93070000",
         129 => x"03474102",
         130 => x"e39407fc",
         131 => x"9307e006",
         132 => x"630af700",
         133 => x"93050000",
         134 => x"13057102",
         135 => x"ef00d001",
         136 => x"13040500",
         137 => x"93773400",
         138 => x"639e0710",
         139 => x"b7170010",
         140 => x"138c87f2",
         141 => x"b7170010",
         142 => x"930c0404",
         143 => x"938bc7f4",
         144 => x"130980ff",
         145 => x"93058000",
         146 => x"13050400",
         147 => x"ef005014",
         148 => x"13050c00",
         149 => x"ef00006e",
         150 => x"83240400",
         151 => x"93058000",
         152 => x"930a8001",
         153 => x"13850400",
         154 => x"ef009012",
         155 => x"13850b00",
         156 => x"ef00406c",
         157 => x"b70d00ff",
         158 => x"33f5b401",
         159 => x"33555501",
         160 => x"3387a900",
         161 => x"03470700",
         162 => x"13777709",
         163 => x"63140700",
         164 => x"1305e002",
         165 => x"938a8aff",
         166 => x"ef00c067",
         167 => x"93dd8d00",
         168 => x"e39c2afd",
         169 => x"13044400",
         170 => x"13050a00",
         171 => x"ef008068",
         172 => x"e31a94f9",
         173 => x"6ff09fec",
         174 => x"b7170010",
         175 => x"138547e3",
         176 => x"ef004067",
         177 => x"e38c04ea",
         178 => x"6ff01ff2",
         179 => x"93050000",
         180 => x"13050000",
         181 => x"ef000061",
         182 => x"b70700f0",
         183 => x"23a20700",
         184 => x"93020000",
         185 => x"73905230",
         186 => x"83278101",
         187 => x"e7800700",
         188 => x"e38604e8",
         189 => x"6ff05fef",
         190 => x"03476102",
         191 => x"93070002",
         192 => x"e314f7ea",
         193 => x"93050000",
         194 => x"13057102",
         195 => x"ef00c072",
         196 => x"93773500",
         197 => x"13040500",
         198 => x"63960702",
         199 => x"93058000",
         200 => x"ef001007",
         201 => x"b7170010",
         202 => x"138587f2",
         203 => x"ef008060",
         204 => x"03250400",
         205 => x"93058000",
         206 => x"ef009005",
         207 => x"e38004e4",
         208 => x"6ff09fea",
         209 => x"b7170010",
         210 => x"1385c7f2",
         211 => x"ef00805e",
         212 => x"e38604e2",
         213 => x"6ff05fe9",
         214 => x"03476102",
         215 => x"93070002",
         216 => x"e31af7e4",
         217 => x"b305e100",
         218 => x"13057102",
         219 => x"ef00c06c",
         220 => x"93773500",
         221 => x"13040500",
         222 => x"e39607fc",
         223 => x"03250102",
         224 => x"93050000",
         225 => x"ef00406b",
         226 => x"2320a400",
         227 => x"e38804de",
         228 => x"6ff09fe5",
         229 => x"b70700f0",
         230 => x"23a20700",
         231 => x"93050000",
         232 => x"ef004054",
         233 => x"e7000400",
         234 => x"6ff09fd6",
         235 => x"93041000",
         236 => x"b71c0010",
         237 => x"93878ce2",
         238 => x"232c0100",
         239 => x"370400f0",
         240 => x"13093005",
         241 => x"930aa004",
         242 => x"130b3002",
         243 => x"9309a000",
         244 => x"2326f100",
         245 => x"83274400",
         246 => x"93c71700",
         247 => x"2322f400",
         248 => x"ef00c034",
         249 => x"9377f50f",
         250 => x"63882703",
         251 => x"63825707",
         252 => x"63806709",
         253 => x"e39004fe",
         254 => x"0325c100",
         255 => x"ef008053",
         256 => x"83274400",
         257 => x"93c71700",
         258 => x"2322f400",
         259 => x"ef000032",
         260 => x"9377f50f",
         261 => x"e39c27fd",
         262 => x"ef004031",
         263 => x"937bf50f",
         264 => x"9387fbfc",
         265 => x"93f7f70f",
         266 => x"13072000",
         267 => x"637af704",
         268 => x"93879bfc",
         269 => x"93f7f70f",
         270 => x"13072000",
         271 => x"6370f710",
         272 => x"ef00c02e",
         273 => x"9377f50f",
         274 => x"e39c37ff",
         275 => x"6ff09ffa",
         276 => x"63820416",
         277 => x"93050000",
         278 => x"13050000",
         279 => x"ef008048",
         280 => x"b70700f0",
         281 => x"23a20700",
         282 => x"83278101",
         283 => x"e7800700",
         284 => x"b70700f0",
         285 => x"1307a00a",
         286 => x"23a2e700",
         287 => x"6ff01fcb",
         288 => x"93071003",
         289 => x"638afb16",
         290 => x"93072003",
         291 => x"13052000",
         292 => x"638efb0e",
         293 => x"ef00004e",
         294 => x"930bb5ff",
         295 => x"13058000",
         296 => x"ef00404d",
         297 => x"130d0500",
         298 => x"338cab01",
         299 => x"63840b12",
         300 => x"b70701ff",
         301 => x"9387f7ff",
         302 => x"b7060001",
         303 => x"232af100",
         304 => x"9387f6ff",
         305 => x"232ef100",
         306 => x"b707ffff",
         307 => x"9387f70f",
         308 => x"2328f100",
         309 => x"930b2000",
         310 => x"6f008003",
         311 => x"93073000",
         312 => x"6300f60e",
         313 => x"83270101",
         314 => x"137807f0",
         315 => x"93158500",
         316 => x"3377f700",
         317 => x"93071000",
         318 => x"33650501",
         319 => x"6314f600",
         320 => x"33e5e500",
         321 => x"23a0ad00",
         322 => x"130d1d00",
         323 => x"63048d0d",
         324 => x"13052000",
         325 => x"ef000046",
         326 => x"937dcdff",
         327 => x"13763d00",
         328 => x"03a70d00",
         329 => x"e31c76fb",
         330 => x"83274101",
         331 => x"13150501",
         332 => x"3377f700",
         333 => x"3365e500",
         334 => x"6ff0dffc",
         335 => x"13050700",
         336 => x"ef004043",
         337 => x"93077003",
         338 => x"6380fb0a",
         339 => x"93078003",
         340 => x"638afb04",
         341 => x"13054000",
         342 => x"ef00c041",
         343 => x"930b0500",
         344 => x"130ca000",
         345 => x"ef00801c",
         346 => x"9377f50f",
         347 => x"e39c87ff",
         348 => x"232c7101",
         349 => x"6ff01fe8",
         350 => x"b71c0010",
         351 => x"13858ce2",
         352 => x"ef00403b",
         353 => x"93040000",
         354 => x"6ff0dfe2",
         355 => x"ef00803e",
         356 => x"930bc5ff",
         357 => x"13056000",
         358 => x"ef00c03d",
         359 => x"130d0500",
         360 => x"6ff09ff0",
         361 => x"13056000",
         362 => x"ef00c03c",
         363 => x"930b0500",
         364 => x"6ff01ffb",
         365 => x"13858ce2",
         366 => x"ef00c037",
         367 => x"6ff09fe9",
         368 => x"8327c101",
         369 => x"13158501",
         370 => x"3377f700",
         371 => x"3365e500",
         372 => x"6ff05ff3",
         373 => x"930ba000",
         374 => x"ef004015",
         375 => x"9377f50f",
         376 => x"e39c77ff",
         377 => x"6ff01fe1",
         378 => x"13058000",
         379 => x"ef008038",
         380 => x"930b0500",
         381 => x"6ff0dff6",
         382 => x"13050700",
         383 => x"ef008037",
         384 => x"930bd5ff",
         385 => x"13054000",
         386 => x"ef00c036",
         387 => x"130d0500",
         388 => x"6ff09fe9",
         389 => x"130101fb",
         390 => x"23261104",
         391 => x"23245104",
         392 => x"23226104",
         393 => x"23207104",
         394 => x"232e8102",
         395 => x"232c9102",
         396 => x"232aa102",
         397 => x"2328b102",
         398 => x"2326c102",
         399 => x"2324d102",
         400 => x"2322e102",
         401 => x"2320f102",
         402 => x"232e0101",
         403 => x"232c1101",
         404 => x"232ac101",
         405 => x"2328d101",
         406 => x"2326e101",
         407 => x"2324f101",
         408 => x"73241034",
         409 => x"f3272034",
         410 => x"37150010",
         411 => x"130505dd",
         412 => x"93840700",
         413 => x"ef00002c",
         414 => x"13850400",
         415 => x"93058000",
         416 => x"ef000051",
         417 => x"37150010",
         418 => x"1305c5d5",
         419 => x"ef00802a",
         420 => x"13044400",
         421 => x"73101434",
         422 => x"0324c103",
         423 => x"8320c104",
         424 => x"83228104",
         425 => x"03234104",
         426 => x"83230104",
         427 => x"83248103",
         428 => x"03254103",
         429 => x"83250103",
         430 => x"0326c102",
         431 => x"83268102",
         432 => x"03274102",
         433 => x"83270102",
         434 => x"0328c101",
         435 => x"83288101",
         436 => x"032e4101",
         437 => x"832e0101",
         438 => x"032fc100",
         439 => x"832f8100",
         440 => x"13010105",
         441 => x"73002030",
         442 => x"6f000000",
         443 => x"13030500",
         444 => x"630a0600",
         445 => x"2300b300",
         446 => x"1306f6ff",
         447 => x"13031300",
         448 => x"e31a06fe",
         449 => x"67800000",
         450 => x"13030500",
         451 => x"630e0600",
         452 => x"83830500",
         453 => x"23007300",
         454 => x"1306f6ff",
         455 => x"13031300",
         456 => x"93851500",
         457 => x"e31606fe",
         458 => x"67800000",
         459 => x"370700f0",
         460 => x"13070710",
         461 => x"83274700",
         462 => x"93f78700",
         463 => x"e38c07fe",
         464 => x"03258700",
         465 => x"1375f50f",
         466 => x"67800000",
         467 => x"130101fd",
         468 => x"23202103",
         469 => x"b7170010",
         470 => x"37190010",
         471 => x"23248102",
         472 => x"23229102",
         473 => x"232e3101",
         474 => x"232c4101",
         475 => x"232a5101",
         476 => x"23286101",
         477 => x"23267101",
         478 => x"23261102",
         479 => x"138bf5ff",
         480 => x"930a0500",
         481 => x"1309c9c0",
         482 => x"938b07d6",
         483 => x"13040000",
         484 => x"93045001",
         485 => x"93092000",
         486 => x"130a2001",
         487 => x"eff01ff9",
         488 => x"93070500",
         489 => x"1375f50f",
         490 => x"63c0a402",
         491 => x"63d2a902",
         492 => x"1307d5ff",
         493 => x"636eea00",
         494 => x"13172700",
         495 => x"3307e900",
         496 => x"03270700",
         497 => x"67000700",
         498 => x"1307f007",
         499 => x"6308e506",
         500 => x"635c640f",
         501 => x"138707fe",
         502 => x"1377f70f",
         503 => x"9306e005",
         504 => x"e3eee6fa",
         505 => x"33878a00",
         506 => x"2300f700",
         507 => x"13041400",
         508 => x"ef004012",
         509 => x"6ff09ffa",
         510 => x"b38a8a00",
         511 => x"37150010",
         512 => x"23800a00",
         513 => x"1305c5d5",
         514 => x"ef00c012",
         515 => x"8320c102",
         516 => x"13050400",
         517 => x"03248102",
         518 => x"83244102",
         519 => x"03290102",
         520 => x"8329c101",
         521 => x"032a8101",
         522 => x"832a4101",
         523 => x"032b0101",
         524 => x"832bc100",
         525 => x"13010103",
         526 => x"67800000",
         527 => x"63528006",
         528 => x"1305f007",
         529 => x"ef00000d",
         530 => x"1304f4ff",
         531 => x"6ff01ff5",
         532 => x"13850b00",
         533 => x"ef00000e",
         534 => x"eff05fed",
         535 => x"93070500",
         536 => x"1375f50f",
         537 => x"63c8a402",
         538 => x"13040000",
         539 => x"6ff01ff4",
         540 => x"635c8002",
         541 => x"1305f007",
         542 => x"1304f4ff",
         543 => x"ef008009",
         544 => x"e31a04fe",
         545 => x"eff09fea",
         546 => x"93070500",
         547 => x"1375f50f",
         548 => x"e3dca4fc",
         549 => x"1307f007",
         550 => x"13040000",
         551 => x"e31ae5f2",
         552 => x"13057000",
         553 => x"ef000007",
         554 => x"eff05fe8",
         555 => x"93070500",
         556 => x"13075001",
         557 => x"1375f50f",
         558 => x"e35aa7ee",
         559 => x"1307f007",
         560 => x"e300e5fe",
         561 => x"e34864f1",
         562 => x"13057000",
         563 => x"ef008004",
         564 => x"6ff0dfec",
         565 => x"b70700f0",
         566 => x"03a54710",
         567 => x"13758500",
         568 => x"67800000",
         569 => x"f32710fc",
         570 => x"63960700",
         571 => x"b7f7fa02",
         572 => x"93870708",
         573 => x"63060500",
         574 => x"33d5a702",
         575 => x"1305f5ff",
         576 => x"b70700f0",
         577 => x"23a6a710",
         578 => x"23a0b710",
         579 => x"23a20710",
         580 => x"67800000",
         581 => x"370700f0",
         582 => x"1375f50f",
         583 => x"13070710",
         584 => x"2324a700",
         585 => x"83274700",
         586 => x"93f70701",
         587 => x"e38c07fe",
         588 => x"67800000",
         589 => x"630e0502",
         590 => x"130101ff",
         591 => x"23248100",
         592 => x"23261100",
         593 => x"13040500",
         594 => x"03450500",
         595 => x"630a0500",
         596 => x"13041400",
         597 => x"eff01ffc",
         598 => x"03450400",
         599 => x"e31a05fe",
         600 => x"8320c100",
         601 => x"03248100",
         602 => x"13010101",
         603 => x"67800000",
         604 => x"67800000",
         605 => x"130101fe",
         606 => x"232e1100",
         607 => x"232c8100",
         608 => x"6350a00a",
         609 => x"23263101",
         610 => x"b7190010",
         611 => x"232a9100",
         612 => x"23282101",
         613 => x"23244101",
         614 => x"13090500",
         615 => x"938999c5",
         616 => x"93040000",
         617 => x"13040000",
         618 => x"130a1000",
         619 => x"6f000001",
         620 => x"3364c400",
         621 => x"93841400",
         622 => x"63029904",
         623 => x"eff01fd7",
         624 => x"b387a900",
         625 => x"83c70700",
         626 => x"130605fd",
         627 => x"13144400",
         628 => x"13f74700",
         629 => x"93f64704",
         630 => x"e31c07fc",
         631 => x"93f73700",
         632 => x"e38a06fc",
         633 => x"63944701",
         634 => x"13050502",
         635 => x"130595fa",
         636 => x"93841400",
         637 => x"3364a400",
         638 => x"e31299fc",
         639 => x"8320c101",
         640 => x"13050400",
         641 => x"03248101",
         642 => x"83244101",
         643 => x"03290101",
         644 => x"8329c100",
         645 => x"032a8100",
         646 => x"13010102",
         647 => x"67800000",
         648 => x"13040000",
         649 => x"8320c101",
         650 => x"13050400",
         651 => x"03248101",
         652 => x"13010102",
         653 => x"67800000",
         654 => x"83470500",
         655 => x"37160010",
         656 => x"130696c5",
         657 => x"3307f600",
         658 => x"03470700",
         659 => x"93060500",
         660 => x"13758700",
         661 => x"630e0500",
         662 => x"83c71600",
         663 => x"93861600",
         664 => x"3307f600",
         665 => x"03470700",
         666 => x"13758700",
         667 => x"e31605fe",
         668 => x"13754704",
         669 => x"63040506",
         670 => x"13050000",
         671 => x"13031000",
         672 => x"6f000002",
         673 => x"83c71600",
         674 => x"93861600",
         675 => x"33e5a800",
         676 => x"3307f600",
         677 => x"03470700",
         678 => x"13784704",
         679 => x"63000804",
         680 => x"13784700",
         681 => x"938807fd",
         682 => x"13773700",
         683 => x"13154500",
         684 => x"e31a08fc",
         685 => x"63146700",
         686 => x"93870702",
         687 => x"938797fa",
         688 => x"93861600",
         689 => x"33e5a700",
         690 => x"83c70600",
         691 => x"3307f600",
         692 => x"03470700",
         693 => x"13784704",
         694 => x"e31408fc",
         695 => x"63840500",
         696 => x"23a0d500",
         697 => x"67800000",
         698 => x"130101fd",
         699 => x"23261102",
         700 => x"232a0100",
         701 => x"232c0100",
         702 => x"232e0100",
         703 => x"63000508",
         704 => x"93070500",
         705 => x"63400506",
         706 => x"b7d5cccc",
         707 => x"13850700",
         708 => x"9385d5cc",
         709 => x"93064101",
         710 => x"93089000",
         711 => x"b337b502",
         712 => x"13060500",
         713 => x"13880600",
         714 => x"9386f6ff",
         715 => x"93d73700",
         716 => x"13972700",
         717 => x"3307f700",
         718 => x"13171700",
         719 => x"3305e540",
         720 => x"13050503",
         721 => x"a385a600",
         722 => x"13850700",
         723 => x"e3e8c8fc",
         724 => x"1305a800",
         725 => x"eff01fde",
         726 => x"8320c102",
         727 => x"13010103",
         728 => x"67800000",
         729 => x"2326a100",
         730 => x"1305d002",
         731 => x"eff09fda",
         732 => x"8327c100",
         733 => x"b307f040",
         734 => x"6ff01ff9",
         735 => x"13050003",
         736 => x"eff05fd9",
         737 => x"8320c102",
         738 => x"13010103",
         739 => x"67800000",
         740 => x"130101fe",
         741 => x"232e1100",
         742 => x"23220100",
         743 => x"23240100",
         744 => x"23060100",
         745 => x"1387f5ff",
         746 => x"93077000",
         747 => x"93060500",
         748 => x"63e4e704",
         749 => x"93070700",
         750 => x"13054100",
         751 => x"b307f500",
         752 => x"b385b740",
         753 => x"13089003",
         754 => x"13f6f600",
         755 => x"13070603",
         756 => x"6374e800",
         757 => x"13077605",
         758 => x"2380e700",
         759 => x"9387f7ff",
         760 => x"93d64600",
         761 => x"e392f5fe",
         762 => x"eff0dfd4",
         763 => x"8320c101",
         764 => x"13010102",
         765 => x"67800000",
         766 => x"93058000",
         767 => x"6ff0dffb",
         768 => x"37150010",
         769 => x"1305c5d6",
         770 => x"6ff0dfd2",
         771 => x"50080010",
         772 => x"d0070010",
         773 => x"d0070010",
         774 => x"d0070010",
         775 => x"d0070010",
         776 => x"3c080010",
         777 => x"d0070010",
         778 => x"f8070010",
         779 => x"d0070010",
         780 => x"d0070010",
         781 => x"f8070010",
         782 => x"d0070010",
         783 => x"d0070010",
         784 => x"d0070010",
         785 => x"d0070010",
         786 => x"d0070010",
         787 => x"d0070010",
         788 => x"d0070010",
         789 => x"70080010",
         790 => x"00202020",
         791 => x"20202020",
         792 => x"20202828",
         793 => x"28282820",
         794 => x"20202020",
         795 => x"20202020",
         796 => x"20202020",
         797 => x"20202020",
         798 => x"20881010",
         799 => x"10101010",
         800 => x"10101010",
         801 => x"10101010",
         802 => x"10040404",
         803 => x"04040404",
         804 => x"04040410",
         805 => x"10101010",
         806 => x"10104141",
         807 => x"41414141",
         808 => x"01010101",
         809 => x"01010101",
         810 => x"01010101",
         811 => x"01010101",
         812 => x"01010101",
         813 => x"10101010",
         814 => x"10104242",
         815 => x"42424242",
         816 => x"02020202",
         817 => x"02020202",
         818 => x"02020202",
         819 => x"02020202",
         820 => x"02020202",
         821 => x"10101010",
         822 => x"20000000",
         823 => x"00000000",
         824 => x"00000000",
         825 => x"00000000",
         826 => x"00000000",
         827 => x"00000000",
         828 => x"00000000",
         829 => x"00000000",
         830 => x"00000000",
         831 => x"00000000",
         832 => x"00000000",
         833 => x"00000000",
         834 => x"00000000",
         835 => x"00000000",
         836 => x"00000000",
         837 => x"00000000",
         838 => x"00000000",
         839 => x"00000000",
         840 => x"00000000",
         841 => x"00000000",
         842 => x"00000000",
         843 => x"00000000",
         844 => x"00000000",
         845 => x"00000000",
         846 => x"00000000",
         847 => x"00000000",
         848 => x"00000000",
         849 => x"00000000",
         850 => x"00000000",
         851 => x"00000000",
         852 => x"00000000",
         853 => x"00000000",
         854 => x"00000000",
         855 => x"0d0a0000",
         856 => x"3c627265",
         857 => x"616b3e0d",
         858 => x"0a000000",
         859 => x"0d0a5f5f",
         860 => x"5f202020",
         861 => x"20202020",
         862 => x"5f20205f",
         863 => x"5f202020",
         864 => x"205f205c",
         865 => x"202f5f5f",
         866 => x"205f5f20",
         867 => x"0d0a207c",
         868 => x"207c5f7c",
         869 => x"7c207c7c",
         870 => x"5f7c285f",
         871 => x"202d2d2d",
         872 => x"7c5f2920",
         873 => x"56205f5f",
         874 => x"29205f29",
         875 => x"0d0a207c",
         876 => x"207c207c",
         877 => x"7c5f7c7c",
         878 => x"207c5f5f",
         879 => x"29202020",
         880 => x"7c205c20",
         881 => x"20205f5f",
         882 => x"292f5f5f",
         883 => x"0d0a0000",
         884 => x"54726170",
         885 => x"3a206d63",
         886 => x"61757365",
         887 => x"203d2030",
         888 => x"78000000",
         889 => x"0d0a5448",
         890 => x"55415320",
         891 => x"52495343",
         892 => x"2d562042",
         893 => x"6f6f746c",
         894 => x"6f616465",
         895 => x"72207630",
         896 => x"2e362e34",
         897 => x"0d0a4861",
         898 => x"72647761",
         899 => x"72653a20",
         900 => x"00000000",
         901 => x"0d0a436c",
         902 => x"6f636b20",
         903 => x"66726571",
         904 => x"75656e63",
         905 => x"793a2000",
         906 => x"3f0a0000",
         907 => x"3e200000",
         908 => x"68000000",
         909 => x"48656c70",
         910 => x"3a0d0a20",
         911 => x"68202020",
         912 => x"20202020",
         913 => x"20202020",
         914 => x"20202020",
         915 => x"202d2074",
         916 => x"68697320",
         917 => x"68656c70",
         918 => x"0d0a2072",
         919 => x"20202020",
         920 => x"20202020",
         921 => x"20202020",
         922 => x"20202020",
         923 => x"2d207275",
         924 => x"6e206170",
         925 => x"706c6963",
         926 => x"6174696f",
         927 => x"6e0d0a20",
         928 => x"7277203c",
         929 => x"61646472",
         930 => x"3e202020",
         931 => x"20202020",
         932 => x"202d2072",
         933 => x"65616420",
         934 => x"776f7264",
         935 => x"2066726f",
         936 => x"6d206164",
         937 => x"64720d0a",
         938 => x"20777720",
         939 => x"3c616464",
         940 => x"723e203c",
         941 => x"64617461",
         942 => x"3e202d20",
         943 => x"77726974",
         944 => x"6520776f",
         945 => x"72642064",
         946 => x"61746120",
         947 => x"61742061",
         948 => x"6464720d",
         949 => x"0a206477",
         950 => x"203c6164",
         951 => x"64723e20",
         952 => x"20202020",
         953 => x"2020202d",
         954 => x"2064756d",
         955 => x"70203136",
         956 => x"20776f72",
         957 => x"64730d0a",
         958 => x"206e2020",
         959 => x"20202020",
         960 => x"20202020",
         961 => x"20202020",
         962 => x"20202d20",
         963 => x"64756d70",
         964 => x"206e6578",
         965 => x"74203136",
         966 => x"20776f72",
         967 => x"64730000",
         968 => x"72000000",
         969 => x"72772000",
         970 => x"3a200000",
         971 => x"4e6f7420",
         972 => x"6f6e2034",
         973 => x"2d627974",
         974 => x"6520626f",
         975 => x"756e6461",
         976 => x"72792100",
         977 => x"77772000",
         978 => x"64772000",
         979 => x"20200000",
         980 => x"3f3f0000"
            );
end package bootrom_image;
