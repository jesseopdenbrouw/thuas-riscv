-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Thu Apr 18 10:26:21 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382022f",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"13868187",
           8 => x"9387819e",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13858187",
          13 => x"ef00806c",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93878187",
          17 => x"637cf600",
          18 => x"b7450000",
          19 => x"3386c740",
          20 => x"938545f1",
          21 => x"13050500",
          22 => x"ef00006c",
          23 => x"ef20005a",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef00d029",
          29 => x"ef101045",
          30 => x"6f00901e",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef009022",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"232c4101",
          40 => x"130a0500",
          41 => x"37450000",
          42 => x"130505c6",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"13044100",
          50 => x"ef005020",
          51 => x"37490000",
          52 => x"9309c1ff",
          53 => x"93070400",
          54 => x"130949ae",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef00d01c",
          65 => x"37450000",
          66 => x"130545c7",
          67 => x"ef00101c",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef009019",
          78 => x"37450000",
          79 => x"130505c8",
          80 => x"ef00d018",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74708",
          91 => x"b70600f0",
          92 => x"1377f7fe",
          93 => x"23a2e708",
          94 => x"83a74600",
          95 => x"93c71700",
          96 => x"23a2f600",
          97 => x"67800000",
          98 => x"370700f0",
          99 => x"83274700",
         100 => x"93e70720",
         101 => x"2322f700",
         102 => x"6f000000",
         103 => x"b70700f0",
         104 => x"b70500f0",
         105 => x"370500f0",
         106 => x"9387470f",
         107 => x"9385050f",
         108 => x"83a60700",
         109 => x"03a60500",
         110 => x"03a70700",
         111 => x"e31ad7fe",
         112 => x"b7870100",
         113 => x"b70500f0",
         114 => x"1308f0ff",
         115 => x"9387076a",
         116 => x"23ae050f",
         117 => x"b307f600",
         118 => x"b70600f0",
         119 => x"23ac060f",
         120 => x"33b6c700",
         121 => x"23acf60e",
         122 => x"3306e600",
         123 => x"23aec50e",
         124 => x"83274500",
         125 => x"93c72700",
         126 => x"2322f500",
         127 => x"67800000",
         128 => x"b70700f0",
         129 => x"03a74702",
         130 => x"b70600f0",
         131 => x"93870702",
         132 => x"13778700",
         133 => x"630a0700",
         134 => x"03a74600",
         135 => x"13478700",
         136 => x"23a2e600",
         137 => x"83a78700",
         138 => x"67800000",
         139 => x"b70700f0",
         140 => x"03a7470a",
         141 => x"b70600f0",
         142 => x"1377f7f0",
         143 => x"23a2e70a",
         144 => x"83a74600",
         145 => x"93c74700",
         146 => x"23a2f600",
         147 => x"67800000",
         148 => x"b70700f0",
         149 => x"03a74706",
         150 => x"b70600f0",
         151 => x"137777ff",
         152 => x"23a2e706",
         153 => x"83a74600",
         154 => x"93c70701",
         155 => x"23a2f600",
         156 => x"67800000",
         157 => x"b70700f0",
         158 => x"03a74704",
         159 => x"b70600f0",
         160 => x"137777ff",
         161 => x"23a2e704",
         162 => x"83a74600",
         163 => x"93c70702",
         164 => x"23a2f600",
         165 => x"67800000",
         166 => x"b70700f0",
         167 => x"03a74705",
         168 => x"b70600f0",
         169 => x"137777ff",
         170 => x"23aae704",
         171 => x"83a74600",
         172 => x"93c70708",
         173 => x"23a2f600",
         174 => x"67800000",
         175 => x"b70700f0",
         176 => x"23ae0700",
         177 => x"03a74700",
         178 => x"13470704",
         179 => x"23a2e700",
         180 => x"67800000",
         181 => x"370700f0",
         182 => x"b70600f0",
         183 => x"2326070e",
         184 => x"83a74600",
         185 => x"93c70710",
         186 => x"23a2f600",
         187 => x"67800000",
         188 => x"6f000000",
         189 => x"13050000",
         190 => x"67800000",
         191 => x"13050000",
         192 => x"67800000",
         193 => x"130101f7",
         194 => x"23221100",
         195 => x"23242100",
         196 => x"23263100",
         197 => x"23284100",
         198 => x"232a5100",
         199 => x"232c6100",
         200 => x"232e7100",
         201 => x"23208102",
         202 => x"23229102",
         203 => x"2324a102",
         204 => x"2326b102",
         205 => x"2328c102",
         206 => x"232ad102",
         207 => x"232ce102",
         208 => x"232ef102",
         209 => x"23200105",
         210 => x"23221105",
         211 => x"23242105",
         212 => x"23263105",
         213 => x"23284105",
         214 => x"232a5105",
         215 => x"232c6105",
         216 => x"232e7105",
         217 => x"23208107",
         218 => x"23229107",
         219 => x"2324a107",
         220 => x"2326b107",
         221 => x"2328c107",
         222 => x"232ad107",
         223 => x"232ce107",
         224 => x"232ef107",
         225 => x"f3222034",
         226 => x"23205108",
         227 => x"f3221034",
         228 => x"23225108",
         229 => x"83a20200",
         230 => x"23245108",
         231 => x"f3223034",
         232 => x"23265108",
         233 => x"f3272034",
         234 => x"1307b000",
         235 => x"6374f70c",
         236 => x"37070080",
         237 => x"1307d7ff",
         238 => x"b387e700",
         239 => x"13078001",
         240 => x"636ef700",
         241 => x"37470000",
         242 => x"93972700",
         243 => x"130787af",
         244 => x"b387e700",
         245 => x"83a70700",
         246 => x"67800700",
         247 => x"03258102",
         248 => x"83220108",
         249 => x"63c80200",
         250 => x"f3221034",
         251 => x"93824200",
         252 => x"73901234",
         253 => x"832fc107",
         254 => x"032f8107",
         255 => x"832e4107",
         256 => x"032e0107",
         257 => x"832dc106",
         258 => x"032d8106",
         259 => x"832c4106",
         260 => x"032c0106",
         261 => x"832bc105",
         262 => x"032b8105",
         263 => x"832a4105",
         264 => x"032a0105",
         265 => x"8329c104",
         266 => x"03298104",
         267 => x"83284104",
         268 => x"03280104",
         269 => x"8327c103",
         270 => x"03278103",
         271 => x"83264103",
         272 => x"03260103",
         273 => x"8325c102",
         274 => x"83244102",
         275 => x"03240102",
         276 => x"8323c101",
         277 => x"03238101",
         278 => x"83224101",
         279 => x"03220101",
         280 => x"8321c100",
         281 => x"03218100",
         282 => x"83204100",
         283 => x"13010109",
         284 => x"73002030",
         285 => x"93061000",
         286 => x"e3f2f6f6",
         287 => x"e360f7f6",
         288 => x"37470000",
         289 => x"93972700",
         290 => x"1307c7b5",
         291 => x"b387e700",
         292 => x"83a70700",
         293 => x"67800700",
         294 => x"eff09fdb",
         295 => x"03258102",
         296 => x"6ff01ff4",
         297 => x"eff01fe3",
         298 => x"03258102",
         299 => x"6ff05ff3",
         300 => x"eff0dfce",
         301 => x"03258102",
         302 => x"6ff09ff2",
         303 => x"eff01fe0",
         304 => x"03258102",
         305 => x"6ff0dff1",
         306 => x"eff0dfc9",
         307 => x"03258102",
         308 => x"6ff01ff1",
         309 => x"eff09fd5",
         310 => x"03258102",
         311 => x"6ff05ff0",
         312 => x"eff01fd2",
         313 => x"03258102",
         314 => x"6ff09fef",
         315 => x"eff0dfda",
         316 => x"03258102",
         317 => x"6ff0dfee",
         318 => x"eff0dfd7",
         319 => x"03258102",
         320 => x"6ff01fee",
         321 => x"13050100",
         322 => x"eff01fb9",
         323 => x"03258102",
         324 => x"6ff01fed",
         325 => x"9307900a",
         326 => x"6380f814",
         327 => x"63d81703",
         328 => x"9307600d",
         329 => x"638ef818",
         330 => x"938808c0",
         331 => x"9307f000",
         332 => x"63e01705",
         333 => x"b7470000",
         334 => x"9387c7b8",
         335 => x"93982800",
         336 => x"b388f800",
         337 => x"83a70800",
         338 => x"67800700",
         339 => x"938878fc",
         340 => x"93074002",
         341 => x"63ee1701",
         342 => x"b7470000",
         343 => x"9387c7bc",
         344 => x"93982800",
         345 => x"b388f800",
         346 => x"83a70800",
         347 => x"67800700",
         348 => x"ef204008",
         349 => x"93078005",
         350 => x"2320f500",
         351 => x"9307f0ff",
         352 => x"13850700",
         353 => x"6ff0dfe5",
         354 => x"b7270000",
         355 => x"23a2f500",
         356 => x"93070000",
         357 => x"13850700",
         358 => x"6ff09fe4",
         359 => x"93070000",
         360 => x"13850700",
         361 => x"6ff0dfe3",
         362 => x"ef20c004",
         363 => x"93079000",
         364 => x"2320f500",
         365 => x"9307f0ff",
         366 => x"13850700",
         367 => x"6ff05fe2",
         368 => x"ef204003",
         369 => x"9307f001",
         370 => x"2320f500",
         371 => x"9307f0ff",
         372 => x"13850700",
         373 => x"6ff0dfe0",
         374 => x"ef20c001",
         375 => x"9307d000",
         376 => x"2320f500",
         377 => x"9307f0ff",
         378 => x"13850700",
         379 => x"6ff05fdf",
         380 => x"ef204000",
         381 => x"93072000",
         382 => x"2320f500",
         383 => x"9307f0ff",
         384 => x"13850700",
         385 => x"6ff0dfdd",
         386 => x"13090600",
         387 => x"13840500",
         388 => x"635cc000",
         389 => x"b384c500",
         390 => x"eff01fa6",
         391 => x"2300a400",
         392 => x"13041400",
         393 => x"e39a84fe",
         394 => x"13050900",
         395 => x"6ff05fdb",
         396 => x"13090600",
         397 => x"13840500",
         398 => x"e358c0fe",
         399 => x"b384c500",
         400 => x"03450400",
         401 => x"13041400",
         402 => x"eff05fa3",
         403 => x"e39a84fe",
         404 => x"13050900",
         405 => x"6ff0dfd8",
         406 => x"13090000",
         407 => x"93040500",
         408 => x"13040900",
         409 => x"93090900",
         410 => x"93070900",
         411 => x"732410c8",
         412 => x"f32910c0",
         413 => x"f32710c8",
         414 => x"e31af4fe",
         415 => x"37460f00",
         416 => x"13060624",
         417 => x"93060000",
         418 => x"13850900",
         419 => x"93050400",
         420 => x"ef10401c",
         421 => x"37460f00",
         422 => x"23a4a400",
         423 => x"13060624",
         424 => x"93060000",
         425 => x"13850900",
         426 => x"93050400",
         427 => x"ef00904f",
         428 => x"23a0a400",
         429 => x"23a2b400",
         430 => x"13050900",
         431 => x"6ff05fd2",
         432 => x"63180500",
         433 => x"1385819e",
         434 => x"13050500",
         435 => x"6ff05fd1",
         436 => x"b7870020",
         437 => x"93870700",
         438 => x"13070040",
         439 => x"b387e740",
         440 => x"e364f5fe",
         441 => x"ef101071",
         442 => x"9307c000",
         443 => x"2320f500",
         444 => x"1305f0ff",
         445 => x"13050500",
         446 => x"6ff09fce",
         447 => x"13030500",
         448 => x"630a0600",
         449 => x"2300b300",
         450 => x"1306f6ff",
         451 => x"13031300",
         452 => x"e31a06fe",
         453 => x"67800000",
         454 => x"13030500",
         455 => x"630e0600",
         456 => x"83830500",
         457 => x"23007300",
         458 => x"1306f6ff",
         459 => x"13031300",
         460 => x"93851500",
         461 => x"e31606fe",
         462 => x"67800000",
         463 => x"630c0602",
         464 => x"13030500",
         465 => x"93061000",
         466 => x"636ab500",
         467 => x"9306f0ff",
         468 => x"1307f6ff",
         469 => x"3303e300",
         470 => x"b385e500",
         471 => x"83830500",
         472 => x"23007300",
         473 => x"1306f6ff",
         474 => x"3303d300",
         475 => x"b385d500",
         476 => x"e31606fe",
         477 => x"67800000",
         478 => x"6f000000",
         479 => x"130101ff",
         480 => x"23248100",
         481 => x"13040000",
         482 => x"23229100",
         483 => x"23202101",
         484 => x"23261100",
         485 => x"93040500",
         486 => x"13090400",
         487 => x"93070400",
         488 => x"732410c8",
         489 => x"732910c0",
         490 => x"f32710c8",
         491 => x"e31af4fe",
         492 => x"37460f00",
         493 => x"13060624",
         494 => x"93060000",
         495 => x"13050900",
         496 => x"93050400",
         497 => x"ef100009",
         498 => x"37460f00",
         499 => x"23a4a400",
         500 => x"93050400",
         501 => x"13050900",
         502 => x"13060624",
         503 => x"93060000",
         504 => x"ef00503c",
         505 => x"8320c100",
         506 => x"03248100",
         507 => x"23a0a400",
         508 => x"23a2b400",
         509 => x"03290100",
         510 => x"83244100",
         511 => x"13050000",
         512 => x"13010101",
         513 => x"67800000",
         514 => x"13050000",
         515 => x"67800000",
         516 => x"13050000",
         517 => x"67800000",
         518 => x"130101ff",
         519 => x"23202101",
         520 => x"23261100",
         521 => x"13090600",
         522 => x"6356c002",
         523 => x"23248100",
         524 => x"23229100",
         525 => x"13840500",
         526 => x"b384c500",
         527 => x"03450400",
         528 => x"13041400",
         529 => x"eff09f83",
         530 => x"e39a84fe",
         531 => x"03248100",
         532 => x"83244100",
         533 => x"8320c100",
         534 => x"13050900",
         535 => x"03290100",
         536 => x"13010101",
         537 => x"67800000",
         538 => x"130101ff",
         539 => x"23202101",
         540 => x"23261100",
         541 => x"13090600",
         542 => x"6356c002",
         543 => x"23248100",
         544 => x"23229100",
         545 => x"13840500",
         546 => x"b384c500",
         547 => x"eff0cffe",
         548 => x"13041400",
         549 => x"a30fa4fe",
         550 => x"e39a84fe",
         551 => x"03248100",
         552 => x"83244100",
         553 => x"8320c100",
         554 => x"13050900",
         555 => x"03290100",
         556 => x"13010101",
         557 => x"67800000",
         558 => x"13051000",
         559 => x"67800000",
         560 => x"130101ff",
         561 => x"23261100",
         562 => x"ef10d052",
         563 => x"8320c100",
         564 => x"93076001",
         565 => x"2320f500",
         566 => x"1305f0ff",
         567 => x"13010101",
         568 => x"67800000",
         569 => x"1305f0ff",
         570 => x"67800000",
         571 => x"b7270000",
         572 => x"23a2f500",
         573 => x"13050000",
         574 => x"67800000",
         575 => x"13051000",
         576 => x"67800000",
         577 => x"13050000",
         578 => x"67800000",
         579 => x"130101fe",
         580 => x"2324c100",
         581 => x"2326d100",
         582 => x"2328e100",
         583 => x"232af100",
         584 => x"232c0101",
         585 => x"232e1101",
         586 => x"1305f0ff",
         587 => x"13010102",
         588 => x"67800000",
         589 => x"130101ff",
         590 => x"23261100",
         591 => x"ef10904b",
         592 => x"8320c100",
         593 => x"9307a000",
         594 => x"2320f500",
         595 => x"1305f0ff",
         596 => x"13010101",
         597 => x"67800000",
         598 => x"130101ff",
         599 => x"23261100",
         600 => x"ef105049",
         601 => x"8320c100",
         602 => x"93072000",
         603 => x"2320f500",
         604 => x"1305f0ff",
         605 => x"13010101",
         606 => x"67800000",
         607 => x"b7270000",
         608 => x"23a2f500",
         609 => x"13050000",
         610 => x"67800000",
         611 => x"130101ff",
         612 => x"23261100",
         613 => x"ef101046",
         614 => x"8320c100",
         615 => x"9307f001",
         616 => x"2320f500",
         617 => x"1305f0ff",
         618 => x"13010101",
         619 => x"67800000",
         620 => x"130101ff",
         621 => x"23261100",
         622 => x"ef10d043",
         623 => x"8320c100",
         624 => x"9307b000",
         625 => x"2320f500",
         626 => x"1305f0ff",
         627 => x"13010101",
         628 => x"67800000",
         629 => x"130101ff",
         630 => x"23261100",
         631 => x"ef109041",
         632 => x"8320c100",
         633 => x"9307c000",
         634 => x"2320f500",
         635 => x"1305f0ff",
         636 => x"13010101",
         637 => x"67800000",
         638 => x"03a7c187",
         639 => x"b7870020",
         640 => x"93870700",
         641 => x"93060040",
         642 => x"b387d740",
         643 => x"630c0700",
         644 => x"3305a700",
         645 => x"63e2a702",
         646 => x"23aea186",
         647 => x"13050700",
         648 => x"67800000",
         649 => x"9386819e",
         650 => x"1387819e",
         651 => x"23aed186",
         652 => x"3305a700",
         653 => x"e3f2a7fe",
         654 => x"130101ff",
         655 => x"23261100",
         656 => x"ef10503b",
         657 => x"8320c100",
         658 => x"9307c000",
         659 => x"2320f500",
         660 => x"1307f0ff",
         661 => x"13050700",
         662 => x"13010101",
         663 => x"67800000",
         664 => x"370700f0",
         665 => x"13070702",
         666 => x"83274700",
         667 => x"93f78700",
         668 => x"e38c07fe",
         669 => x"03258700",
         670 => x"1375f50f",
         671 => x"67800000",
         672 => x"f32710fc",
         673 => x"63960700",
         674 => x"b7f7fa02",
         675 => x"93870708",
         676 => x"63060500",
         677 => x"33d5a702",
         678 => x"1305f5ff",
         679 => x"b70700f0",
         680 => x"23a6a702",
         681 => x"23a0b702",
         682 => x"67800000",
         683 => x"370700f0",
         684 => x"1375f50f",
         685 => x"13070702",
         686 => x"2324a700",
         687 => x"83274700",
         688 => x"93f70701",
         689 => x"e38c07fe",
         690 => x"67800000",
         691 => x"630e0502",
         692 => x"130101ff",
         693 => x"23248100",
         694 => x"23261100",
         695 => x"13040500",
         696 => x"03450500",
         697 => x"630a0500",
         698 => x"13041400",
         699 => x"eff01ffc",
         700 => x"03450400",
         701 => x"e31a05fe",
         702 => x"8320c100",
         703 => x"03248100",
         704 => x"13010101",
         705 => x"67800000",
         706 => x"67800000",
         707 => x"130101f9",
         708 => x"23229106",
         709 => x"23202107",
         710 => x"23261106",
         711 => x"23248106",
         712 => x"232e3105",
         713 => x"232c4105",
         714 => x"232a5105",
         715 => x"23286105",
         716 => x"23267105",
         717 => x"23248105",
         718 => x"23229105",
         719 => x"2320a105",
         720 => x"13090500",
         721 => x"93840500",
         722 => x"232c0100",
         723 => x"232e0100",
         724 => x"23200102",
         725 => x"23220102",
         726 => x"23240102",
         727 => x"23260102",
         728 => x"23280102",
         729 => x"232a0102",
         730 => x"232c0102",
         731 => x"232e0102",
         732 => x"732410fc",
         733 => x"63160400",
         734 => x"37f4fa02",
         735 => x"13040408",
         736 => x"97f2ffff",
         737 => x"93824278",
         738 => x"73905230",
         739 => x"37c50100",
         740 => x"93059000",
         741 => x"13050520",
         742 => x"eff09fee",
         743 => x"b7270000",
         744 => x"93870771",
         745 => x"b356f402",
         746 => x"13561400",
         747 => x"370700f0",
         748 => x"1306f6ff",
         749 => x"b7170300",
         750 => x"2326c708",
         751 => x"130e1001",
         752 => x"938707d4",
         753 => x"2320c709",
         754 => x"370600f0",
         755 => x"37230000",
         756 => x"1303f370",
         757 => x"37581200",
         758 => x"130808f8",
         759 => x"b70800f0",
         760 => x"370500f0",
         761 => x"b70500f0",
         762 => x"3357f402",
         763 => x"9387f6ff",
         764 => x"2328f60a",
         765 => x"2326660a",
         766 => x"2320c60b",
         767 => x"93078070",
         768 => x"23a0f806",
         769 => x"b3570403",
         770 => x"1307f7ff",
         771 => x"13170701",
         772 => x"13678700",
         773 => x"2320e504",
         774 => x"1307a007",
         775 => x"9387f7ff",
         776 => x"93970701",
         777 => x"93e7c700",
         778 => x"23a8f504",
         779 => x"b70700f0",
         780 => x"23ace700",
         781 => x"f3224030",
         782 => x"93e20208",
         783 => x"73904230",
         784 => x"f3224030",
         785 => x"93e28200",
         786 => x"73904230",
         787 => x"b7220000",
         788 => x"93828280",
         789 => x"73900230",
         790 => x"b7490000",
         791 => x"138509c8",
         792 => x"eff0dfe6",
         793 => x"1304f9ff",
         794 => x"63522003",
         795 => x"1309f0ff",
         796 => x"03a50400",
         797 => x"1304f4ff",
         798 => x"93844400",
         799 => x"eff01fe5",
         800 => x"138509c8",
         801 => x"eff09fe4",
         802 => x"e31424ff",
         803 => x"37450000",
         804 => x"130545c8",
         805 => x"37f9eeee",
         806 => x"b7faeeee",
         807 => x"b7090010",
         808 => x"37140000",
         809 => x"eff09fe2",
         810 => x"374b0000",
         811 => x"9389f9ff",
         812 => x"1309f9ee",
         813 => x"938aeaee",
         814 => x"130404e1",
         815 => x"93040000",
         816 => x"b71b0000",
         817 => x"938b0b2c",
         818 => x"130af000",
         819 => x"6f00c000",
         820 => x"938bfbff",
         821 => x"63840b18",
         822 => x"93050000",
         823 => x"13058100",
         824 => x"ef10101e",
         825 => x"e31605fe",
         826 => x"032c8100",
         827 => x"8325c100",
         828 => x"13060400",
         829 => x"9357cc01",
         830 => x"13974500",
         831 => x"b367f700",
         832 => x"b3f73701",
         833 => x"33773c01",
         834 => x"13d5f541",
         835 => x"13d88501",
         836 => x"3307f700",
         837 => x"33070701",
         838 => x"9377d500",
         839 => x"3307f700",
         840 => x"33774703",
         841 => x"937725ff",
         842 => x"93860400",
         843 => x"13050c00",
         844 => x"938bfbff",
         845 => x"3307f700",
         846 => x"b307ec40",
         847 => x"1357f741",
         848 => x"3338fc00",
         849 => x"3387e540",
         850 => x"33070741",
         851 => x"b3885703",
         852 => x"33072703",
         853 => x"33b82703",
         854 => x"33071701",
         855 => x"b3872703",
         856 => x"33070701",
         857 => x"1358f741",
         858 => x"13783800",
         859 => x"b307f800",
         860 => x"33b80701",
         861 => x"3307e800",
         862 => x"1318e701",
         863 => x"93d72700",
         864 => x"b367f800",
         865 => x"13582740",
         866 => x"93184800",
         867 => x"13d3c701",
         868 => x"33e36800",
         869 => x"33733301",
         870 => x"b3f83701",
         871 => x"135e8801",
         872 => x"1357f741",
         873 => x"b3886800",
         874 => x"b388c801",
         875 => x"1373d700",
         876 => x"b3886800",
         877 => x"b3f84803",
         878 => x"137727ff",
         879 => x"939c4700",
         880 => x"b38cfc40",
         881 => x"939c2c00",
         882 => x"b30c9c41",
         883 => x"b388e800",
         884 => x"33871741",
         885 => x"93d8f841",
         886 => x"33b3e700",
         887 => x"33081841",
         888 => x"33086840",
         889 => x"33082803",
         890 => x"33035703",
         891 => x"b3382703",
         892 => x"33086800",
         893 => x"33072703",
         894 => x"33081801",
         895 => x"9358f841",
         896 => x"93f83800",
         897 => x"3387e800",
         898 => x"b3381701",
         899 => x"b3880801",
         900 => x"9398e801",
         901 => x"13572700",
         902 => x"33e7e800",
         903 => x"13184700",
         904 => x"3307e840",
         905 => x"13172700",
         906 => x"338de740",
         907 => x"ef00c007",
         908 => x"83260101",
         909 => x"13070500",
         910 => x"13880c00",
         911 => x"93070d00",
         912 => x"13060c00",
         913 => x"93054bcb",
         914 => x"13058101",
         915 => x"ef10c038",
         916 => x"13058101",
         917 => x"eff09fc7",
         918 => x"e3900be8",
         919 => x"73001000",
         920 => x"b70700f0",
         921 => x"9306f00f",
         922 => x"23a4d706",
         923 => x"370700f0",
         924 => x"83260704",
         925 => x"93050009",
         926 => x"b70700f0",
         927 => x"93e60630",
         928 => x"2320d704",
         929 => x"2324b704",
         930 => x"03a60705",
         931 => x"b70600f0",
         932 => x"13660630",
         933 => x"23a8c704",
         934 => x"23acb704",
         935 => x"93071000",
         936 => x"23a6f60e",
         937 => x"6ff0dfe1",
         938 => x"13080000",
         939 => x"63c60512",
         940 => x"63dc0600",
         941 => x"b337c000",
         942 => x"b306d040",
         943 => x"1348f8ff",
         944 => x"b386f640",
         945 => x"3306c040",
         946 => x"93080600",
         947 => x"13070500",
         948 => x"13830500",
         949 => x"639a060e",
         950 => x"63f4c516",
         951 => x"b7070100",
         952 => x"6364f622",
         953 => x"b7070001",
         954 => x"93068001",
         955 => x"6374f600",
         956 => x"93060001",
         957 => x"335ed600",
         958 => x"97370000",
         959 => x"938747ec",
         960 => x"b387c701",
         961 => x"83c70700",
         962 => x"130e0002",
         963 => x"b387d700",
         964 => x"b306fe40",
         965 => x"630cfe00",
         966 => x"3393d500",
         967 => x"b357f500",
         968 => x"b318d600",
         969 => x"33e36700",
         970 => x"3317d500",
         971 => x"13d60801",
         972 => x"3355c302",
         973 => x"93960801",
         974 => x"93d60601",
         975 => x"93570701",
         976 => x"3373c302",
         977 => x"b385a602",
         978 => x"13130301",
         979 => x"b3e76700",
         980 => x"63fcb700",
         981 => x"b387f800",
         982 => x"1303f5ff",
         983 => x"63e41701",
         984 => x"63e6b742",
         985 => x"13050300",
         986 => x"b387b740",
         987 => x"b3d5c702",
         988 => x"13170701",
         989 => x"13570701",
         990 => x"b3f7c702",
         991 => x"b386b602",
         992 => x"93970701",
         993 => x"3367f700",
         994 => x"637ed700",
         995 => x"3387e800",
         996 => x"9387f5ff",
         997 => x"63661701",
         998 => x"9385e5ff",
         999 => x"6364d700",
        1000 => x"93850700",
        1001 => x"13150501",
        1002 => x"3365b500",
        1003 => x"93050000",
        1004 => x"630a0800",
        1005 => x"b337a000",
        1006 => x"b305b040",
        1007 => x"b385f540",
        1008 => x"3305a040",
        1009 => x"67800000",
        1010 => x"63f4d502",
        1011 => x"93050000",
        1012 => x"13050000",
        1013 => x"6ff0dffd",
        1014 => x"b337a000",
        1015 => x"b305b040",
        1016 => x"b385f540",
        1017 => x"3305a040",
        1018 => x"1308f0ff",
        1019 => x"6ff05fec",
        1020 => x"b7070100",
        1021 => x"63e8f61e",
        1022 => x"37070001",
        1023 => x"93078001",
        1024 => x"63f4e600",
        1025 => x"93070001",
        1026 => x"b3d8f600",
        1027 => x"17370000",
        1028 => x"130707db",
        1029 => x"33071701",
        1030 => x"03470700",
        1031 => x"13030002",
        1032 => x"3307f700",
        1033 => x"b308e340",
        1034 => x"6316e31e",
        1035 => x"63e4b632",
        1036 => x"3335c500",
        1037 => x"13351500",
        1038 => x"93050000",
        1039 => x"6ff05ff7",
        1040 => x"630c060c",
        1041 => x"b7070100",
        1042 => x"637cf62e",
        1043 => x"13330610",
        1044 => x"13331300",
        1045 => x"13133300",
        1046 => x"b3566600",
        1047 => x"97370000",
        1048 => x"938707d6",
        1049 => x"b387d700",
        1050 => x"83c60700",
        1051 => x"93070002",
        1052 => x"b3866600",
        1053 => x"b38ed740",
        1054 => x"6394d70c",
        1055 => x"b386c540",
        1056 => x"13530601",
        1057 => x"13160601",
        1058 => x"13560601",
        1059 => x"93051000",
        1060 => x"33d56602",
        1061 => x"93570701",
        1062 => x"b3f66602",
        1063 => x"330ec502",
        1064 => x"93960601",
        1065 => x"b3e7d700",
        1066 => x"63fcc701",
        1067 => x"b387f800",
        1068 => x"9306f5ff",
        1069 => x"63e41701",
        1070 => x"63e4c72d",
        1071 => x"13850600",
        1072 => x"b387c741",
        1073 => x"b3d66702",
        1074 => x"13170701",
        1075 => x"13570701",
        1076 => x"b3f76702",
        1077 => x"3386c602",
        1078 => x"93970701",
        1079 => x"3367f700",
        1080 => x"637ec700",
        1081 => x"3387e800",
        1082 => x"9387f6ff",
        1083 => x"63661701",
        1084 => x"9386e6ff",
        1085 => x"6364c700",
        1086 => x"93860700",
        1087 => x"13150501",
        1088 => x"3365d500",
        1089 => x"6ff0dfea",
        1090 => x"93360610",
        1091 => x"93b61600",
        1092 => x"93963600",
        1093 => x"6ff01fde",
        1094 => x"93060000",
        1095 => x"97370000",
        1096 => x"938707ca",
        1097 => x"b387d700",
        1098 => x"83c60700",
        1099 => x"13030000",
        1100 => x"93070002",
        1101 => x"b3866600",
        1102 => x"b38ed740",
        1103 => x"e380d7f4",
        1104 => x"b318d601",
        1105 => x"33ded500",
        1106 => x"13d30801",
        1107 => x"b3576e02",
        1108 => x"13960801",
        1109 => x"13560601",
        1110 => x"b356d500",
        1111 => x"3317d501",
        1112 => x"b395d501",
        1113 => x"b3e6b600",
        1114 => x"93d50601",
        1115 => x"337e6e02",
        1116 => x"3305f602",
        1117 => x"131e0e01",
        1118 => x"b3e5c501",
        1119 => x"63fea500",
        1120 => x"b385b800",
        1121 => x"138ef7ff",
        1122 => x"63e4151f",
        1123 => x"63f2a51e",
        1124 => x"9387e7ff",
        1125 => x"b3851501",
        1126 => x"b385a540",
        1127 => x"33d56502",
        1128 => x"93960601",
        1129 => x"93d60601",
        1130 => x"b3f56502",
        1131 => x"330ea602",
        1132 => x"93950501",
        1133 => x"b3e6b600",
        1134 => x"63fec601",
        1135 => x"b386d800",
        1136 => x"9305f5ff",
        1137 => x"63ee1619",
        1138 => x"63fcc619",
        1139 => x"1305e5ff",
        1140 => x"b3861601",
        1141 => x"93950701",
        1142 => x"b386c641",
        1143 => x"b3e5a500",
        1144 => x"6ff01feb",
        1145 => x"93b70610",
        1146 => x"93b71700",
        1147 => x"93973700",
        1148 => x"b3d8f600",
        1149 => x"17370000",
        1150 => x"130787bc",
        1151 => x"33071701",
        1152 => x"03470700",
        1153 => x"13030002",
        1154 => x"3307f700",
        1155 => x"b308e340",
        1156 => x"e30ee3e0",
        1157 => x"b35ee600",
        1158 => x"b3961601",
        1159 => x"b3eede00",
        1160 => x"33d3e500",
        1161 => x"13df0e01",
        1162 => x"b357e303",
        1163 => x"139e0e01",
        1164 => x"b3951501",
        1165 => x"135e0e01",
        1166 => x"3357e500",
        1167 => x"3367b700",
        1168 => x"93560701",
        1169 => x"33161601",
        1170 => x"3373e303",
        1171 => x"b305fe02",
        1172 => x"13130301",
        1173 => x"b3e66600",
        1174 => x"63feb600",
        1175 => x"b386de00",
        1176 => x"1383f7ff",
        1177 => x"63ead611",
        1178 => x"63f8b610",
        1179 => x"9387e7ff",
        1180 => x"b386d601",
        1181 => x"b386b640",
        1182 => x"b3d5e603",
        1183 => x"13170701",
        1184 => x"13570701",
        1185 => x"b3f6e603",
        1186 => x"3303be02",
        1187 => x"93960601",
        1188 => x"3367d700",
        1189 => x"637e6700",
        1190 => x"3387ee00",
        1191 => x"9386f5ff",
        1192 => x"6364d70d",
        1193 => x"6372670c",
        1194 => x"9385e5ff",
        1195 => x"3307d701",
        1196 => x"93970701",
        1197 => x"370f0100",
        1198 => x"b3e7b700",
        1199 => x"9306ffff",
        1200 => x"b3f5d700",
        1201 => x"13de0701",
        1202 => x"b376d600",
        1203 => x"13560601",
        1204 => x"b38ed502",
        1205 => x"33076740",
        1206 => x"b306de02",
        1207 => x"13d30e01",
        1208 => x"b385c502",
        1209 => x"b385d500",
        1210 => x"b305b300",
        1211 => x"330ece02",
        1212 => x"63f4d500",
        1213 => x"330eee01",
        1214 => x"93d60501",
        1215 => x"b386c601",
        1216 => x"636ad702",
        1217 => x"6308d700",
        1218 => x"13850700",
        1219 => x"93050000",
        1220 => x"6ff01fca",
        1221 => x"b7060100",
        1222 => x"9386f6ff",
        1223 => x"33f7d500",
        1224 => x"13170701",
        1225 => x"b3fede00",
        1226 => x"33151501",
        1227 => x"3307d701",
        1228 => x"e37ce5fc",
        1229 => x"1385f7ff",
        1230 => x"93050000",
        1231 => x"6ff05fc7",
        1232 => x"b7070001",
        1233 => x"637af604",
        1234 => x"93560601",
        1235 => x"13030001",
        1236 => x"6ff0dfd0",
        1237 => x"93050000",
        1238 => x"13051000",
        1239 => x"6ff05fc5",
        1240 => x"13850500",
        1241 => x"6ff01fe7",
        1242 => x"93850600",
        1243 => x"6ff05ff4",
        1244 => x"93070e00",
        1245 => x"6ff05fe2",
        1246 => x"93070300",
        1247 => x"6ff09fef",
        1248 => x"1305e5ff",
        1249 => x"b3871701",
        1250 => x"6ff09fd3",
        1251 => x"1305e5ff",
        1252 => x"b3871701",
        1253 => x"6ff05fbd",
        1254 => x"93568601",
        1255 => x"13038001",
        1256 => x"6ff0dfcb",
        1257 => x"13080600",
        1258 => x"93080500",
        1259 => x"13870500",
        1260 => x"6390060e",
        1261 => x"63fec512",
        1262 => x"b7070100",
        1263 => x"636ef61e",
        1264 => x"b7070001",
        1265 => x"93068001",
        1266 => x"6374f600",
        1267 => x"93060001",
        1268 => x"3353d600",
        1269 => x"97370000",
        1270 => x"9387879e",
        1271 => x"b3876700",
        1272 => x"83c70700",
        1273 => x"13030002",
        1274 => x"b387d700",
        1275 => x"b306f340",
        1276 => x"630cf300",
        1277 => x"3397d500",
        1278 => x"b357f500",
        1279 => x"3318d600",
        1280 => x"33e7e700",
        1281 => x"b318d500",
        1282 => x"13560801",
        1283 => x"3355c702",
        1284 => x"93160801",
        1285 => x"93d60601",
        1286 => x"93d70801",
        1287 => x"3377c702",
        1288 => x"b385a602",
        1289 => x"13170701",
        1290 => x"b3e7e700",
        1291 => x"63fcb700",
        1292 => x"b307f800",
        1293 => x"1307f5ff",
        1294 => x"63e40701",
        1295 => x"63e0b740",
        1296 => x"13050700",
        1297 => x"b387b740",
        1298 => x"33d7c702",
        1299 => x"93980801",
        1300 => x"93d80801",
        1301 => x"b3f7c702",
        1302 => x"b386e602",
        1303 => x"93970701",
        1304 => x"b3e8f800",
        1305 => x"63fed800",
        1306 => x"b3081801",
        1307 => x"9307f7ff",
        1308 => x"63e60801",
        1309 => x"1307e7ff",
        1310 => x"63e4d800",
        1311 => x"13870700",
        1312 => x"13150501",
        1313 => x"3365e500",
        1314 => x"93050000",
        1315 => x"67800000",
        1316 => x"63f8d500",
        1317 => x"93050000",
        1318 => x"13050000",
        1319 => x"67800000",
        1320 => x"b7070100",
        1321 => x"63e8f61e",
        1322 => x"37070001",
        1323 => x"93078001",
        1324 => x"63f4e600",
        1325 => x"93070001",
        1326 => x"33d8f600",
        1327 => x"17370000",
        1328 => x"13070790",
        1329 => x"33070701",
        1330 => x"03470700",
        1331 => x"93080002",
        1332 => x"3307f700",
        1333 => x"3388e840",
        1334 => x"6396e81e",
        1335 => x"63e4b632",
        1336 => x"3335c500",
        1337 => x"13351500",
        1338 => x"93050000",
        1339 => x"67800000",
        1340 => x"630c060c",
        1341 => x"b7070100",
        1342 => x"637cf62e",
        1343 => x"13370610",
        1344 => x"13371700",
        1345 => x"13173700",
        1346 => x"b356e600",
        1347 => x"97370000",
        1348 => x"9387078b",
        1349 => x"b387d700",
        1350 => x"83c70700",
        1351 => x"93060002",
        1352 => x"b387e700",
        1353 => x"b38ef640",
        1354 => x"6394f60c",
        1355 => x"b387c540",
        1356 => x"93560601",
        1357 => x"13160601",
        1358 => x"13560601",
        1359 => x"93051000",
        1360 => x"33d5d702",
        1361 => x"13d70801",
        1362 => x"b3f7d702",
        1363 => x"3303c502",
        1364 => x"93970701",
        1365 => x"b367f700",
        1366 => x"63fc6700",
        1367 => x"b307f800",
        1368 => x"1307f5ff",
        1369 => x"63e40701",
        1370 => x"63e4672c",
        1371 => x"13050700",
        1372 => x"b3876740",
        1373 => x"33d7d702",
        1374 => x"93980801",
        1375 => x"93d80801",
        1376 => x"b3f7d702",
        1377 => x"3306c702",
        1378 => x"93970701",
        1379 => x"b3e8f800",
        1380 => x"63fec800",
        1381 => x"b3081801",
        1382 => x"9307f7ff",
        1383 => x"63e60801",
        1384 => x"1307e7ff",
        1385 => x"63e4c800",
        1386 => x"13870700",
        1387 => x"13150501",
        1388 => x"3365e500",
        1389 => x"67800000",
        1390 => x"93360610",
        1391 => x"93b61600",
        1392 => x"93963600",
        1393 => x"6ff0dfe0",
        1394 => x"93060000",
        1395 => x"97270000",
        1396 => x"9387077f",
        1397 => x"b387d700",
        1398 => x"83c70700",
        1399 => x"13070000",
        1400 => x"93060002",
        1401 => x"b387e700",
        1402 => x"b38ef640",
        1403 => x"e380f6f4",
        1404 => x"3318d601",
        1405 => x"33d3f500",
        1406 => x"93560801",
        1407 => x"335ed302",
        1408 => x"13160801",
        1409 => x"b395d501",
        1410 => x"13560601",
        1411 => x"b357f500",
        1412 => x"b3e7b700",
        1413 => x"13d70701",
        1414 => x"b318d501",
        1415 => x"3373d302",
        1416 => x"b305c603",
        1417 => x"13130301",
        1418 => x"33676700",
        1419 => x"637eb700",
        1420 => x"3307e800",
        1421 => x"1305feff",
        1422 => x"6364071f",
        1423 => x"6372b71e",
        1424 => x"130eeeff",
        1425 => x"33070701",
        1426 => x"3307b740",
        1427 => x"3355d702",
        1428 => x"93970701",
        1429 => x"93d70701",
        1430 => x"3377d702",
        1431 => x"3303a602",
        1432 => x"13170701",
        1433 => x"b3e7e700",
        1434 => x"63fe6700",
        1435 => x"b307f800",
        1436 => x"1307f5ff",
        1437 => x"63ee0719",
        1438 => x"63fc6718",
        1439 => x"1305e5ff",
        1440 => x"b3870701",
        1441 => x"93150e01",
        1442 => x"b3876740",
        1443 => x"b3e5a500",
        1444 => x"6ff01feb",
        1445 => x"93b70610",
        1446 => x"93b71700",
        1447 => x"93973700",
        1448 => x"33d8f600",
        1449 => x"17270000",
        1450 => x"13078771",
        1451 => x"33070701",
        1452 => x"03470700",
        1453 => x"93080002",
        1454 => x"3307f700",
        1455 => x"3388e840",
        1456 => x"e38ee8e0",
        1457 => x"335ee600",
        1458 => x"b3960601",
        1459 => x"336ede00",
        1460 => x"b3d8e500",
        1461 => x"935e0e01",
        1462 => x"b3d7d803",
        1463 => x"13130e01",
        1464 => x"b3950501",
        1465 => x"13530301",
        1466 => x"3357e500",
        1467 => x"3367b700",
        1468 => x"93560701",
        1469 => x"33160601",
        1470 => x"b3f8d803",
        1471 => x"b305f302",
        1472 => x"93980801",
        1473 => x"b3e61601",
        1474 => x"63feb600",
        1475 => x"b306de00",
        1476 => x"9388f7ff",
        1477 => x"63eac611",
        1478 => x"63f8b610",
        1479 => x"9387e7ff",
        1480 => x"b386c601",
        1481 => x"b386b640",
        1482 => x"b3d5d603",
        1483 => x"13170701",
        1484 => x"13570701",
        1485 => x"b3f6d603",
        1486 => x"b308b302",
        1487 => x"93960601",
        1488 => x"3367d700",
        1489 => x"637e1701",
        1490 => x"3307ee00",
        1491 => x"9386f5ff",
        1492 => x"6364c70d",
        1493 => x"6372170d",
        1494 => x"9385e5ff",
        1495 => x"3307c701",
        1496 => x"93970701",
        1497 => x"b70e0100",
        1498 => x"b3e7b700",
        1499 => x"9386feff",
        1500 => x"b3f5d700",
        1501 => x"13d30701",
        1502 => x"b376d600",
        1503 => x"13560601",
        1504 => x"338ed502",
        1505 => x"33071741",
        1506 => x"b306d302",
        1507 => x"93580e01",
        1508 => x"b385c502",
        1509 => x"b385d500",
        1510 => x"b385b800",
        1511 => x"3303c302",
        1512 => x"63f4d500",
        1513 => x"3303d301",
        1514 => x"93d60501",
        1515 => x"b3866600",
        1516 => x"636ad702",
        1517 => x"6308d700",
        1518 => x"13850700",
        1519 => x"93050000",
        1520 => x"67800000",
        1521 => x"b7060100",
        1522 => x"9386f6ff",
        1523 => x"33f7d500",
        1524 => x"13170701",
        1525 => x"337ede00",
        1526 => x"33150501",
        1527 => x"3307c701",
        1528 => x"e37ce5fc",
        1529 => x"1385f7ff",
        1530 => x"93050000",
        1531 => x"67800000",
        1532 => x"b7070001",
        1533 => x"637af604",
        1534 => x"93560601",
        1535 => x"13070001",
        1536 => x"6ff0dfd0",
        1537 => x"93050000",
        1538 => x"13051000",
        1539 => x"67800000",
        1540 => x"13050700",
        1541 => x"6ff01fe7",
        1542 => x"93850600",
        1543 => x"6ff05ff4",
        1544 => x"130e0500",
        1545 => x"6ff05fe2",
        1546 => x"93870800",
        1547 => x"6ff09fef",
        1548 => x"1305e5ff",
        1549 => x"b3870701",
        1550 => x"6ff09fd3",
        1551 => x"1305e5ff",
        1552 => x"b3870701",
        1553 => x"6ff01fc0",
        1554 => x"93568601",
        1555 => x"13078001",
        1556 => x"6ff0dfcb",
        1557 => x"13080600",
        1558 => x"93080500",
        1559 => x"93870500",
        1560 => x"13870500",
        1561 => x"6398060c",
        1562 => x"63fac512",
        1563 => x"b7070100",
        1564 => x"636cf61c",
        1565 => x"b7070001",
        1566 => x"93068001",
        1567 => x"6374f600",
        1568 => x"93060001",
        1569 => x"3353d600",
        1570 => x"97270000",
        1571 => x"93874753",
        1572 => x"b3876700",
        1573 => x"83c70700",
        1574 => x"13030002",
        1575 => x"b387d700",
        1576 => x"b306f340",
        1577 => x"630cf300",
        1578 => x"3397d500",
        1579 => x"b357f500",
        1580 => x"3318d600",
        1581 => x"33e7e700",
        1582 => x"b318d500",
        1583 => x"93550801",
        1584 => x"3356b702",
        1585 => x"13130801",
        1586 => x"13530301",
        1587 => x"93d70801",
        1588 => x"3377b702",
        1589 => x"33066602",
        1590 => x"13170701",
        1591 => x"b3e7e700",
        1592 => x"63f8c700",
        1593 => x"b307f800",
        1594 => x"63e40701",
        1595 => x"63e2c73c",
        1596 => x"b387c740",
        1597 => x"33d7b702",
        1598 => x"13950801",
        1599 => x"13550501",
        1600 => x"b3f7b702",
        1601 => x"33076702",
        1602 => x"93970701",
        1603 => x"3365f500",
        1604 => x"637ae500",
        1605 => x"3305a800",
        1606 => x"63660501",
        1607 => x"6374e500",
        1608 => x"33050501",
        1609 => x"3305e540",
        1610 => x"3355d500",
        1611 => x"93050000",
        1612 => x"67800000",
        1613 => x"63f4d500",
        1614 => x"67800000",
        1615 => x"37070100",
        1616 => x"63e6e61c",
        1617 => x"37070001",
        1618 => x"13088001",
        1619 => x"63f4e600",
        1620 => x"13080001",
        1621 => x"33d30601",
        1622 => x"17270000",
        1623 => x"13074746",
        1624 => x"33076700",
        1625 => x"03470700",
        1626 => x"13030002",
        1627 => x"33070701",
        1628 => x"3308e340",
        1629 => x"6314e31c",
        1630 => x"63e4b600",
        1631 => x"636ac500",
        1632 => x"b308c540",
        1633 => x"b386d540",
        1634 => x"b3371501",
        1635 => x"b387f640",
        1636 => x"13850800",
        1637 => x"93850700",
        1638 => x"67800000",
        1639 => x"630e060a",
        1640 => x"b7070100",
        1641 => x"6374f62e",
        1642 => x"13370610",
        1643 => x"13371700",
        1644 => x"13173700",
        1645 => x"b356e600",
        1646 => x"97270000",
        1647 => x"93874740",
        1648 => x"b387d700",
        1649 => x"83c70700",
        1650 => x"13030002",
        1651 => x"b387e700",
        1652 => x"b306f340",
        1653 => x"6316f30a",
        1654 => x"3387c540",
        1655 => x"13530601",
        1656 => x"13160601",
        1657 => x"13560601",
        1658 => x"b3556702",
        1659 => x"93d70801",
        1660 => x"33776702",
        1661 => x"b385c502",
        1662 => x"13170701",
        1663 => x"b3e7e700",
        1664 => x"63fab700",
        1665 => x"b307f800",
        1666 => x"63e60701",
        1667 => x"63f4b700",
        1668 => x"b3870701",
        1669 => x"b387b740",
        1670 => x"33d76702",
        1671 => x"93980801",
        1672 => x"93d80801",
        1673 => x"b3f76702",
        1674 => x"3307c702",
        1675 => x"13950701",
        1676 => x"33e5a800",
        1677 => x"e360e5ee",
        1678 => x"3305e540",
        1679 => x"3355d500",
        1680 => x"93050000",
        1681 => x"67800000",
        1682 => x"93360610",
        1683 => x"93b61600",
        1684 => x"93963600",
        1685 => x"6ff01fe3",
        1686 => x"93060000",
        1687 => x"97270000",
        1688 => x"93870736",
        1689 => x"b387d700",
        1690 => x"83c70700",
        1691 => x"13070000",
        1692 => x"13030002",
        1693 => x"b387e700",
        1694 => x"b306f340",
        1695 => x"e30ef3f4",
        1696 => x"3318d600",
        1697 => x"33def500",
        1698 => x"13530801",
        1699 => x"b35e6e02",
        1700 => x"13160801",
        1701 => x"b395d500",
        1702 => x"3357f500",
        1703 => x"13560601",
        1704 => x"3367b700",
        1705 => x"93570701",
        1706 => x"b318d500",
        1707 => x"337e6e02",
        1708 => x"b385ce02",
        1709 => x"131e0e01",
        1710 => x"b3e7c701",
        1711 => x"63fab700",
        1712 => x"b307f800",
        1713 => x"63e60701",
        1714 => x"63f4b700",
        1715 => x"b3870701",
        1716 => x"b387b740",
        1717 => x"b3d56702",
        1718 => x"13170701",
        1719 => x"13570701",
        1720 => x"b3f76702",
        1721 => x"b385c502",
        1722 => x"93970701",
        1723 => x"3367f700",
        1724 => x"637ab700",
        1725 => x"3307e800",
        1726 => x"63660701",
        1727 => x"6374b700",
        1728 => x"33070701",
        1729 => x"3307b740",
        1730 => x"6ff01fee",
        1731 => x"13b80610",
        1732 => x"13381800",
        1733 => x"13183800",
        1734 => x"33d30601",
        1735 => x"17270000",
        1736 => x"1307072a",
        1737 => x"33076700",
        1738 => x"03470700",
        1739 => x"13030002",
        1740 => x"33070701",
        1741 => x"3308e340",
        1742 => x"e300e3e4",
        1743 => x"b3960601",
        1744 => x"b358e600",
        1745 => x"b3e8d800",
        1746 => x"33dee500",
        1747 => x"13df0801",
        1748 => x"b357ee03",
        1749 => x"939e0801",
        1750 => x"93de0e01",
        1751 => x"b356e500",
        1752 => x"33130501",
        1753 => x"b3950501",
        1754 => x"b3e5b600",
        1755 => x"93d60501",
        1756 => x"33160601",
        1757 => x"337eee03",
        1758 => x"3385fe02",
        1759 => x"131e0e01",
        1760 => x"b3e6c601",
        1761 => x"63fea600",
        1762 => x"b386d800",
        1763 => x"138ef7ff",
        1764 => x"63ec1611",
        1765 => x"63faa610",
        1766 => x"9387e7ff",
        1767 => x"b3861601",
        1768 => x"b386a640",
        1769 => x"33d5e603",
        1770 => x"93950501",
        1771 => x"93d50501",
        1772 => x"b3f6e603",
        1773 => x"b38eae02",
        1774 => x"93960601",
        1775 => x"b3e5d500",
        1776 => x"63fed501",
        1777 => x"b385b800",
        1778 => x"9306f5ff",
        1779 => x"63ea150d",
        1780 => x"63f8d50d",
        1781 => x"1305e5ff",
        1782 => x"b3851501",
        1783 => x"93960701",
        1784 => x"b7020100",
        1785 => x"b3e6a600",
        1786 => x"1385f2ff",
        1787 => x"33fea600",
        1788 => x"935f0601",
        1789 => x"93d60601",
        1790 => x"3375a600",
        1791 => x"330fae02",
        1792 => x"b385d541",
        1793 => x"3385a602",
        1794 => x"93570f01",
        1795 => x"330efe03",
        1796 => x"330eae00",
        1797 => x"b387c701",
        1798 => x"b386f603",
        1799 => x"63f4a700",
        1800 => x"b3865600",
        1801 => x"b70e0100",
        1802 => x"938efeff",
        1803 => x"33f5d701",
        1804 => x"13de0701",
        1805 => x"13150501",
        1806 => x"337fdf01",
        1807 => x"b307de00",
        1808 => x"3305e501",
        1809 => x"63e8f502",
        1810 => x"6384f502",
        1811 => x"3305a340",
        1812 => x"3333a300",
        1813 => x"b385f540",
        1814 => x"b3856540",
        1815 => x"3397e500",
        1816 => x"33550501",
        1817 => x"3365a700",
        1818 => x"b3d50501",
        1819 => x"67800000",
        1820 => x"e37ea3fc",
        1821 => x"3306c540",
        1822 => x"3335c500",
        1823 => x"b3081501",
        1824 => x"b3871741",
        1825 => x"13050600",
        1826 => x"6ff05ffc",
        1827 => x"b7070001",
        1828 => x"6374f602",
        1829 => x"93560601",
        1830 => x"13070001",
        1831 => x"6ff0dfd1",
        1832 => x"13850600",
        1833 => x"6ff09ff3",
        1834 => x"93070e00",
        1835 => x"6ff05fef",
        1836 => x"b3870701",
        1837 => x"6ff0dfc3",
        1838 => x"93568601",
        1839 => x"13078001",
        1840 => x"6ff09fcf",
        1841 => x"130101ff",
        1842 => x"23248100",
        1843 => x"23261100",
        1844 => x"93070000",
        1845 => x"13040500",
        1846 => x"63880700",
        1847 => x"93050000",
        1848 => x"97000000",
        1849 => x"e7000000",
        1850 => x"83a70188",
        1851 => x"63840700",
        1852 => x"e7800700",
        1853 => x"13050400",
        1854 => x"efe01fa8",
        1855 => x"130101ff",
        1856 => x"23248100",
        1857 => x"23261100",
        1858 => x"13040500",
        1859 => x"2316b500",
        1860 => x"2317c500",
        1861 => x"23200500",
        1862 => x"23220500",
        1863 => x"23240500",
        1864 => x"23220506",
        1865 => x"23280500",
        1866 => x"232a0500",
        1867 => x"232c0500",
        1868 => x"13068000",
        1869 => x"93050000",
        1870 => x"1305c505",
        1871 => x"efe01f9c",
        1872 => x"97070000",
        1873 => x"93878750",
        1874 => x"2322f402",
        1875 => x"97070000",
        1876 => x"93874755",
        1877 => x"2324f402",
        1878 => x"97070000",
        1879 => x"9387c75c",
        1880 => x"2326f402",
        1881 => x"97070000",
        1882 => x"93878761",
        1883 => x"2328f402",
        1884 => x"23208402",
        1885 => x"97e7ff1f",
        1886 => x"9387c733",
        1887 => x"630af400",
        1888 => x"93878191",
        1889 => x"6306f400",
        1890 => x"93870198",
        1891 => x"631cf400",
        1892 => x"13058405",
        1893 => x"03248100",
        1894 => x"8320c100",
        1895 => x"13010101",
        1896 => x"6f00500f",
        1897 => x"8320c100",
        1898 => x"03248100",
        1899 => x"13010101",
        1900 => x"67800000",
        1901 => x"13868181",
        1902 => x"97250000",
        1903 => x"9385c5a4",
        1904 => x"17e5ff1f",
        1905 => x"13054526",
        1906 => x"6f00c02f",
        1907 => x"83254500",
        1908 => x"130101ff",
        1909 => x"23248100",
        1910 => x"23261100",
        1911 => x"97e7ff1f",
        1912 => x"9387472d",
        1913 => x"13040500",
        1914 => x"6384f500",
        1915 => x"ef109021",
        1916 => x"83258400",
        1917 => x"93878191",
        1918 => x"6386f500",
        1919 => x"13050400",
        1920 => x"ef105020",
        1921 => x"8325c400",
        1922 => x"93870198",
        1923 => x"638cf500",
        1924 => x"13050400",
        1925 => x"03248100",
        1926 => x"8320c100",
        1927 => x"13010101",
        1928 => x"6f10501e",
        1929 => x"8320c100",
        1930 => x"03248100",
        1931 => x"13010101",
        1932 => x"67800000",
        1933 => x"83a74506",
        1934 => x"93f71700",
        1935 => x"63980702",
        1936 => x"83d7c500",
        1937 => x"93f70720",
        1938 => x"63920702",
        1939 => x"03a58505",
        1940 => x"130101ff",
        1941 => x"23261100",
        1942 => x"ef00d004",
        1943 => x"8320c100",
        1944 => x"13050000",
        1945 => x"13010101",
        1946 => x"67800000",
        1947 => x"13050000",
        1948 => x"67800000",
        1949 => x"83a74506",
        1950 => x"93f71700",
        1951 => x"63980702",
        1952 => x"83d7c500",
        1953 => x"93f70720",
        1954 => x"63920702",
        1955 => x"03a58505",
        1956 => x"130101ff",
        1957 => x"23261100",
        1958 => x"ef005002",
        1959 => x"8320c100",
        1960 => x"13050000",
        1961 => x"13010101",
        1962 => x"67800000",
        1963 => x"13050000",
        1964 => x"67800000",
        1965 => x"130101ff",
        1966 => x"97070000",
        1967 => x"9387c7ef",
        1968 => x"13060000",
        1969 => x"93054000",
        1970 => x"17e5ff1f",
        1971 => x"1305851e",
        1972 => x"23261100",
        1973 => x"23a0f188",
        1974 => x"eff05fe2",
        1975 => x"13061000",
        1976 => x"93059000",
        1977 => x"13858191",
        1978 => x"eff05fe1",
        1979 => x"8320c100",
        1980 => x"13062000",
        1981 => x"93052001",
        1982 => x"13850198",
        1983 => x"13010101",
        1984 => x"6ff0dfdf",
        1985 => x"1385418a",
        1986 => x"6f00c079",
        1987 => x"1385418a",
        1988 => x"6f00c07a",
        1989 => x"130101ff",
        1990 => x"23202101",
        1991 => x"23261100",
        1992 => x"23248100",
        1993 => x"23229100",
        1994 => x"13090500",
        1995 => x"eff09ffd",
        1996 => x"83a70188",
        1997 => x"63940700",
        1998 => x"eff0dff7",
        1999 => x"93848181",
        2000 => x"03a48400",
        2001 => x"83a74400",
        2002 => x"9387f7ff",
        2003 => x"63da0702",
        2004 => x"83a70400",
        2005 => x"6398070c",
        2006 => x"9305c01a",
        2007 => x"13050900",
        2008 => x"ef00500f",
        2009 => x"13040500",
        2010 => x"631c0508",
        2011 => x"23a00400",
        2012 => x"eff0dff9",
        2013 => x"9307c000",
        2014 => x"2320f900",
        2015 => x"6f000006",
        2016 => x"0317c400",
        2017 => x"631a0706",
        2018 => x"b707ffff",
        2019 => x"93871700",
        2020 => x"2326f400",
        2021 => x"13058405",
        2022 => x"23220406",
        2023 => x"ef00806f",
        2024 => x"eff0dff6",
        2025 => x"13068000",
        2026 => x"23200400",
        2027 => x"23240400",
        2028 => x"23220400",
        2029 => x"23280400",
        2030 => x"232a0400",
        2031 => x"232c0400",
        2032 => x"93050000",
        2033 => x"1305c405",
        2034 => x"efe04ff3",
        2035 => x"232a0402",
        2036 => x"232c0402",
        2037 => x"23240404",
        2038 => x"23260404",
        2039 => x"8320c100",
        2040 => x"13050400",
        2041 => x"03248100",
        2042 => x"83244100",
        2043 => x"03290100",
        2044 => x"13010101",
        2045 => x"67800000",
        2046 => x"13048406",
        2047 => x"6ff0dff4",
        2048 => x"93074000",
        2049 => x"23200500",
        2050 => x"2322f500",
        2051 => x"1305c500",
        2052 => x"2324a400",
        2053 => x"1306001a",
        2054 => x"93050000",
        2055 => x"efe00fee",
        2056 => x"23a08400",
        2057 => x"83a40400",
        2058 => x"6ff09ff1",
        2059 => x"130101ff",
        2060 => x"23248100",
        2061 => x"23261100",
        2062 => x"13040500",
        2063 => x"eff09fec",
        2064 => x"83270402",
        2065 => x"638a0700",
        2066 => x"03248100",
        2067 => x"8320c100",
        2068 => x"13010101",
        2069 => x"6ff09feb",
        2070 => x"97070000",
        2071 => x"938747d7",
        2072 => x"2320f402",
        2073 => x"83a70188",
        2074 => x"e39007fe",
        2075 => x"eff09fe4",
        2076 => x"6ff09ffd",
        2077 => x"130101ff",
        2078 => x"23261100",
        2079 => x"eff09fe8",
        2080 => x"8320c100",
        2081 => x"13868181",
        2082 => x"97050000",
        2083 => x"9385c5da",
        2084 => x"13050000",
        2085 => x"13010101",
        2086 => x"6f00c002",
        2087 => x"130101ff",
        2088 => x"13868181",
        2089 => x"97050000",
        2090 => x"938505dd",
        2091 => x"13050000",
        2092 => x"23261100",
        2093 => x"ef000001",
        2094 => x"8320c100",
        2095 => x"13010101",
        2096 => x"6ff0dfe4",
        2097 => x"130101fd",
        2098 => x"23248102",
        2099 => x"23202103",
        2100 => x"232e3101",
        2101 => x"232c4101",
        2102 => x"23286101",
        2103 => x"23267101",
        2104 => x"23261102",
        2105 => x"23229102",
        2106 => x"232a5101",
        2107 => x"93090500",
        2108 => x"138a0500",
        2109 => x"13040600",
        2110 => x"13090000",
        2111 => x"130b1000",
        2112 => x"930bf0ff",
        2113 => x"83248400",
        2114 => x"832a4400",
        2115 => x"938afaff",
        2116 => x"63de0a02",
        2117 => x"03240400",
        2118 => x"e31604fe",
        2119 => x"8320c102",
        2120 => x"03248102",
        2121 => x"83244102",
        2122 => x"8329c101",
        2123 => x"032a8101",
        2124 => x"832a4101",
        2125 => x"032b0101",
        2126 => x"832bc100",
        2127 => x"13050900",
        2128 => x"03290102",
        2129 => x"13010103",
        2130 => x"67800000",
        2131 => x"83d7c400",
        2132 => x"637efb00",
        2133 => x"8397e400",
        2134 => x"638a7701",
        2135 => x"93850400",
        2136 => x"13850900",
        2137 => x"e7000a00",
        2138 => x"3369a900",
        2139 => x"93848406",
        2140 => x"6ff0dff9",
        2141 => x"130101f6",
        2142 => x"232af108",
        2143 => x"b7070080",
        2144 => x"9387f7ff",
        2145 => x"232ef100",
        2146 => x"2328f100",
        2147 => x"b707ffff",
        2148 => x"2326d108",
        2149 => x"2324b100",
        2150 => x"232cb100",
        2151 => x"93878720",
        2152 => x"9306c108",
        2153 => x"93058100",
        2154 => x"232e1106",
        2155 => x"232af100",
        2156 => x"2328e108",
        2157 => x"232c0109",
        2158 => x"232e1109",
        2159 => x"2322d100",
        2160 => x"ef009039",
        2161 => x"83278100",
        2162 => x"23800700",
        2163 => x"8320c107",
        2164 => x"1301010a",
        2165 => x"67800000",
        2166 => x"130101f6",
        2167 => x"232af108",
        2168 => x"b7070080",
        2169 => x"9387f7ff",
        2170 => x"232ef100",
        2171 => x"2328f100",
        2172 => x"b707ffff",
        2173 => x"2324c108",
        2174 => x"2326d108",
        2175 => x"2324a100",
        2176 => x"232ca100",
        2177 => x"93878720",
        2178 => x"93068108",
        2179 => x"13860500",
        2180 => x"03a54187",
        2181 => x"93058100",
        2182 => x"232e1106",
        2183 => x"232af100",
        2184 => x"2328e108",
        2185 => x"232c0109",
        2186 => x"232e1109",
        2187 => x"2322d100",
        2188 => x"ef009032",
        2189 => x"83278100",
        2190 => x"23800700",
        2191 => x"8320c107",
        2192 => x"1301010a",
        2193 => x"67800000",
        2194 => x"130101ff",
        2195 => x"23248100",
        2196 => x"13840500",
        2197 => x"8395e500",
        2198 => x"23261100",
        2199 => x"ef008030",
        2200 => x"63400502",
        2201 => x"83274405",
        2202 => x"b387a700",
        2203 => x"232af404",
        2204 => x"8320c100",
        2205 => x"03248100",
        2206 => x"13010101",
        2207 => x"67800000",
        2208 => x"8357c400",
        2209 => x"37f7ffff",
        2210 => x"1307f7ff",
        2211 => x"b3f7e700",
        2212 => x"2316f400",
        2213 => x"6ff0dffd",
        2214 => x"13050000",
        2215 => x"67800000",
        2216 => x"83d7c500",
        2217 => x"130101fe",
        2218 => x"232c8100",
        2219 => x"232a9100",
        2220 => x"23282101",
        2221 => x"23263101",
        2222 => x"232e1100",
        2223 => x"93f70710",
        2224 => x"93040500",
        2225 => x"13840500",
        2226 => x"13090600",
        2227 => x"93890600",
        2228 => x"638a0700",
        2229 => x"8395e500",
        2230 => x"93062000",
        2231 => x"13060000",
        2232 => x"ef00c023",
        2233 => x"8357c400",
        2234 => x"37f7ffff",
        2235 => x"1307f7ff",
        2236 => x"b3f7e700",
        2237 => x"8315e400",
        2238 => x"2316f400",
        2239 => x"03248101",
        2240 => x"8320c101",
        2241 => x"93860900",
        2242 => x"13060900",
        2243 => x"8329c100",
        2244 => x"03290101",
        2245 => x"13850400",
        2246 => x"83244101",
        2247 => x"13010102",
        2248 => x"6f00c028",
        2249 => x"130101ff",
        2250 => x"23248100",
        2251 => x"13840500",
        2252 => x"8395e500",
        2253 => x"23261100",
        2254 => x"ef00401e",
        2255 => x"1307f0ff",
        2256 => x"8357c400",
        2257 => x"6312e502",
        2258 => x"37f7ffff",
        2259 => x"1307f7ff",
        2260 => x"b3f7e700",
        2261 => x"2316f400",
        2262 => x"8320c100",
        2263 => x"03248100",
        2264 => x"13010101",
        2265 => x"67800000",
        2266 => x"37170000",
        2267 => x"b3e7e700",
        2268 => x"2316f400",
        2269 => x"232aa404",
        2270 => x"6ff01ffe",
        2271 => x"8395e500",
        2272 => x"6f004000",
        2273 => x"130101ff",
        2274 => x"23248100",
        2275 => x"13040500",
        2276 => x"13850500",
        2277 => x"23a20188",
        2278 => x"23261100",
        2279 => x"efe08fd4",
        2280 => x"9307f0ff",
        2281 => x"6318f500",
        2282 => x"83a74188",
        2283 => x"63840700",
        2284 => x"2320f400",
        2285 => x"8320c100",
        2286 => x"03248100",
        2287 => x"13010101",
        2288 => x"67800000",
        2289 => x"83a74187",
        2290 => x"6388a714",
        2291 => x"8327c501",
        2292 => x"130101fe",
        2293 => x"232c8100",
        2294 => x"232e1100",
        2295 => x"232a9100",
        2296 => x"23282101",
        2297 => x"23263101",
        2298 => x"13040500",
        2299 => x"638a0704",
        2300 => x"83a7c700",
        2301 => x"638c0702",
        2302 => x"93040000",
        2303 => x"13090008",
        2304 => x"8327c401",
        2305 => x"83a7c700",
        2306 => x"b3879700",
        2307 => x"83a50700",
        2308 => x"639c050c",
        2309 => x"93844400",
        2310 => x"e39424ff",
        2311 => x"8327c401",
        2312 => x"13050400",
        2313 => x"83a5c700",
        2314 => x"ef00802a",
        2315 => x"8327c401",
        2316 => x"83a50700",
        2317 => x"63860500",
        2318 => x"13050400",
        2319 => x"ef004029",
        2320 => x"83254401",
        2321 => x"63860500",
        2322 => x"13050400",
        2323 => x"ef004028",
        2324 => x"8325c401",
        2325 => x"63860500",
        2326 => x"13050400",
        2327 => x"ef004027",
        2328 => x"83250403",
        2329 => x"63860500",
        2330 => x"13050400",
        2331 => x"ef004026",
        2332 => x"83254403",
        2333 => x"63860500",
        2334 => x"13050400",
        2335 => x"ef004025",
        2336 => x"83258403",
        2337 => x"63860500",
        2338 => x"13050400",
        2339 => x"ef004024",
        2340 => x"83258404",
        2341 => x"63860500",
        2342 => x"13050400",
        2343 => x"ef004023",
        2344 => x"83254404",
        2345 => x"63860500",
        2346 => x"13050400",
        2347 => x"ef004022",
        2348 => x"8325c402",
        2349 => x"63860500",
        2350 => x"13050400",
        2351 => x"ef004021",
        2352 => x"83270402",
        2353 => x"638c0702",
        2354 => x"13050400",
        2355 => x"03248101",
        2356 => x"8320c101",
        2357 => x"83244101",
        2358 => x"03290101",
        2359 => x"8329c100",
        2360 => x"13010102",
        2361 => x"67800700",
        2362 => x"83a90500",
        2363 => x"13050400",
        2364 => x"ef00001e",
        2365 => x"93850900",
        2366 => x"6ff09ff1",
        2367 => x"8320c101",
        2368 => x"03248101",
        2369 => x"83244101",
        2370 => x"03290101",
        2371 => x"8329c100",
        2372 => x"13010102",
        2373 => x"67800000",
        2374 => x"67800000",
        2375 => x"130101ff",
        2376 => x"23248100",
        2377 => x"13040500",
        2378 => x"13850500",
        2379 => x"93050600",
        2380 => x"13860600",
        2381 => x"23a20188",
        2382 => x"23261100",
        2383 => x"efe08fbc",
        2384 => x"9307f0ff",
        2385 => x"6318f500",
        2386 => x"83a74188",
        2387 => x"63840700",
        2388 => x"2320f400",
        2389 => x"8320c100",
        2390 => x"03248100",
        2391 => x"13010101",
        2392 => x"67800000",
        2393 => x"130101ff",
        2394 => x"23248100",
        2395 => x"13040500",
        2396 => x"13850500",
        2397 => x"93050600",
        2398 => x"13860600",
        2399 => x"23a20188",
        2400 => x"23261100",
        2401 => x"efe04fae",
        2402 => x"9307f0ff",
        2403 => x"6318f500",
        2404 => x"83a74188",
        2405 => x"63840700",
        2406 => x"2320f400",
        2407 => x"8320c100",
        2408 => x"03248100",
        2409 => x"13010101",
        2410 => x"67800000",
        2411 => x"130101ff",
        2412 => x"23248100",
        2413 => x"13040500",
        2414 => x"13850500",
        2415 => x"93050600",
        2416 => x"13860600",
        2417 => x"23a20188",
        2418 => x"23261100",
        2419 => x"efe0cfa4",
        2420 => x"9307f0ff",
        2421 => x"6318f500",
        2422 => x"83a74188",
        2423 => x"63840700",
        2424 => x"2320f400",
        2425 => x"8320c100",
        2426 => x"03248100",
        2427 => x"13010101",
        2428 => x"67800000",
        2429 => x"03a54187",
        2430 => x"67800000",
        2431 => x"130101ff",
        2432 => x"23248100",
        2433 => x"23229100",
        2434 => x"17240000",
        2435 => x"1304c490",
        2436 => x"97240000",
        2437 => x"93844490",
        2438 => x"b3848440",
        2439 => x"23202101",
        2440 => x"23261100",
        2441 => x"93d42440",
        2442 => x"13090000",
        2443 => x"631e9902",
        2444 => x"17240000",
        2445 => x"1304448e",
        2446 => x"97240000",
        2447 => x"9384c48d",
        2448 => x"b3848440",
        2449 => x"93d42440",
        2450 => x"13090000",
        2451 => x"63189902",
        2452 => x"8320c100",
        2453 => x"03248100",
        2454 => x"83244100",
        2455 => x"03290100",
        2456 => x"13010101",
        2457 => x"67800000",
        2458 => x"83270400",
        2459 => x"13091900",
        2460 => x"13044400",
        2461 => x"e7800700",
        2462 => x"6ff05ffb",
        2463 => x"83270400",
        2464 => x"13091900",
        2465 => x"13044400",
        2466 => x"e7800700",
        2467 => x"6ff01ffc",
        2468 => x"67800000",
        2469 => x"67800000",
        2470 => x"67800000",
        2471 => x"67800000",
        2472 => x"67800000",
        2473 => x"67800000",
        2474 => x"13051000",
        2475 => x"67800000",
        2476 => x"13051000",
        2477 => x"67800000",
        2478 => x"67800000",
        2479 => x"67800000",
        2480 => x"13860500",
        2481 => x"93050500",
        2482 => x"03a54187",
        2483 => x"6f108022",
        2484 => x"638c050e",
        2485 => x"83a7c5ff",
        2486 => x"130101fe",
        2487 => x"232c8100",
        2488 => x"232e1100",
        2489 => x"1384c5ff",
        2490 => x"63d40700",
        2491 => x"3304f400",
        2492 => x"2326a100",
        2493 => x"ef004032",
        2494 => x"1387c18a",
        2495 => x"83270700",
        2496 => x"0325c100",
        2497 => x"639e0700",
        2498 => x"23220400",
        2499 => x"23208700",
        2500 => x"03248101",
        2501 => x"8320c101",
        2502 => x"13010102",
        2503 => x"6f004030",
        2504 => x"6374f402",
        2505 => x"03260400",
        2506 => x"b306c400",
        2507 => x"639ad700",
        2508 => x"83a60700",
        2509 => x"83a74700",
        2510 => x"b386c600",
        2511 => x"2320d400",
        2512 => x"2322f400",
        2513 => x"6ff09ffc",
        2514 => x"13870700",
        2515 => x"83a74700",
        2516 => x"63840700",
        2517 => x"e37af4fe",
        2518 => x"83260700",
        2519 => x"3306d700",
        2520 => x"63188602",
        2521 => x"03260400",
        2522 => x"b386c600",
        2523 => x"2320d700",
        2524 => x"3306d700",
        2525 => x"e39ec7f8",
        2526 => x"03a60700",
        2527 => x"83a74700",
        2528 => x"b306d600",
        2529 => x"2320d700",
        2530 => x"2322f700",
        2531 => x"6ff05ff8",
        2532 => x"6378c400",
        2533 => x"9307c000",
        2534 => x"2320f500",
        2535 => x"6ff05ff7",
        2536 => x"03260400",
        2537 => x"b306c400",
        2538 => x"639ad700",
        2539 => x"83a60700",
        2540 => x"83a74700",
        2541 => x"b386c600",
        2542 => x"2320d400",
        2543 => x"2322f400",
        2544 => x"23228700",
        2545 => x"6ff0dff4",
        2546 => x"67800000",
        2547 => x"130101ff",
        2548 => x"23202101",
        2549 => x"1389818a",
        2550 => x"83270900",
        2551 => x"23248100",
        2552 => x"23229100",
        2553 => x"23261100",
        2554 => x"93040500",
        2555 => x"13840500",
        2556 => x"63980700",
        2557 => x"93050000",
        2558 => x"ef100014",
        2559 => x"2320a900",
        2560 => x"93050400",
        2561 => x"13850400",
        2562 => x"ef100013",
        2563 => x"1309f0ff",
        2564 => x"63122503",
        2565 => x"1304f0ff",
        2566 => x"8320c100",
        2567 => x"13050400",
        2568 => x"03248100",
        2569 => x"83244100",
        2570 => x"03290100",
        2571 => x"13010101",
        2572 => x"67800000",
        2573 => x"13043500",
        2574 => x"1374c4ff",
        2575 => x"e30e85fc",
        2576 => x"b305a440",
        2577 => x"13850400",
        2578 => x"ef10000f",
        2579 => x"e31625fd",
        2580 => x"6ff05ffc",
        2581 => x"130101fe",
        2582 => x"232a9100",
        2583 => x"93843500",
        2584 => x"93f4c4ff",
        2585 => x"23282101",
        2586 => x"232e1100",
        2587 => x"232c8100",
        2588 => x"23263101",
        2589 => x"23244101",
        2590 => x"93848400",
        2591 => x"9307c000",
        2592 => x"13090500",
        2593 => x"63f2f40a",
        2594 => x"9304c000",
        2595 => x"63e0b40a",
        2596 => x"13050900",
        2597 => x"ef004018",
        2598 => x"9389c18a",
        2599 => x"83a70900",
        2600 => x"13840700",
        2601 => x"631a040a",
        2602 => x"93850400",
        2603 => x"13050900",
        2604 => x"eff0dff1",
        2605 => x"9307f0ff",
        2606 => x"13040500",
        2607 => x"6316f514",
        2608 => x"03a40900",
        2609 => x"93070400",
        2610 => x"639c0710",
        2611 => x"63040412",
        2612 => x"032a0400",
        2613 => x"93050000",
        2614 => x"13050900",
        2615 => x"330a4401",
        2616 => x"ef108005",
        2617 => x"6318aa10",
        2618 => x"83270400",
        2619 => x"13050900",
        2620 => x"b384f440",
        2621 => x"93850400",
        2622 => x"eff05fed",
        2623 => x"9307f0ff",
        2624 => x"630af50e",
        2625 => x"83270400",
        2626 => x"b3879700",
        2627 => x"2320f400",
        2628 => x"83a70900",
        2629 => x"638e070e",
        2630 => x"03a74700",
        2631 => x"6318870c",
        2632 => x"23a20700",
        2633 => x"6f004006",
        2634 => x"e3d204f6",
        2635 => x"9307c000",
        2636 => x"2320f900",
        2637 => x"13050000",
        2638 => x"8320c101",
        2639 => x"03248101",
        2640 => x"83244101",
        2641 => x"03290101",
        2642 => x"8329c100",
        2643 => x"032a8100",
        2644 => x"13010102",
        2645 => x"67800000",
        2646 => x"83260400",
        2647 => x"b3869640",
        2648 => x"63ca0606",
        2649 => x"1307b000",
        2650 => x"637ad704",
        2651 => x"23209400",
        2652 => x"33079400",
        2653 => x"63908704",
        2654 => x"23a0e900",
        2655 => x"83274400",
        2656 => x"2320d700",
        2657 => x"2322f700",
        2658 => x"13050900",
        2659 => x"ef004009",
        2660 => x"1305b400",
        2661 => x"93074400",
        2662 => x"137585ff",
        2663 => x"3307f540",
        2664 => x"e30cf5f8",
        2665 => x"3304e400",
        2666 => x"b387a740",
        2667 => x"2320f400",
        2668 => x"6ff09ff8",
        2669 => x"23a2e700",
        2670 => x"6ff05ffc",
        2671 => x"03274400",
        2672 => x"63968700",
        2673 => x"23a0e900",
        2674 => x"6ff01ffc",
        2675 => x"23a2e700",
        2676 => x"6ff09ffb",
        2677 => x"93070400",
        2678 => x"03244400",
        2679 => x"6ff09fec",
        2680 => x"13840700",
        2681 => x"83a74700",
        2682 => x"6ff01fee",
        2683 => x"93070700",
        2684 => x"6ff05ff2",
        2685 => x"9307c000",
        2686 => x"2320f900",
        2687 => x"13050900",
        2688 => x"ef000002",
        2689 => x"6ff01ff3",
        2690 => x"23209500",
        2691 => x"6ff0dff7",
        2692 => x"23220000",
        2693 => x"73001000",
        2694 => x"13858189",
        2695 => x"6ff09fc8",
        2696 => x"13858189",
        2697 => x"6ff09fc9",
        2698 => x"130101fe",
        2699 => x"23282101",
        2700 => x"03a98500",
        2701 => x"232c8100",
        2702 => x"23263101",
        2703 => x"23225101",
        2704 => x"23206101",
        2705 => x"232e1100",
        2706 => x"232a9100",
        2707 => x"23244101",
        2708 => x"83aa0500",
        2709 => x"13840500",
        2710 => x"130b0600",
        2711 => x"93890600",
        2712 => x"63ec2609",
        2713 => x"8397c500",
        2714 => x"13f70748",
        2715 => x"63040708",
        2716 => x"03274401",
        2717 => x"93043000",
        2718 => x"83a50501",
        2719 => x"b384e402",
        2720 => x"13072000",
        2721 => x"b38aba40",
        2722 => x"130a0500",
        2723 => x"b3c4e402",
        2724 => x"13871600",
        2725 => x"33075701",
        2726 => x"63f4e400",
        2727 => x"93040700",
        2728 => x"93f70740",
        2729 => x"6386070a",
        2730 => x"93850400",
        2731 => x"13050a00",
        2732 => x"eff05fda",
        2733 => x"13090500",
        2734 => x"630c050a",
        2735 => x"83250401",
        2736 => x"13860a00",
        2737 => x"efd05fc5",
        2738 => x"8357c400",
        2739 => x"93f7f7b7",
        2740 => x"93e70708",
        2741 => x"2316f400",
        2742 => x"23282401",
        2743 => x"232a9400",
        2744 => x"33095901",
        2745 => x"b3845441",
        2746 => x"23202401",
        2747 => x"23249400",
        2748 => x"13890900",
        2749 => x"63f42901",
        2750 => x"13890900",
        2751 => x"03250400",
        2752 => x"13060900",
        2753 => x"93050b00",
        2754 => x"efd05fc3",
        2755 => x"83278400",
        2756 => x"13050000",
        2757 => x"b3872741",
        2758 => x"2324f400",
        2759 => x"83270400",
        2760 => x"b3872701",
        2761 => x"2320f400",
        2762 => x"8320c101",
        2763 => x"03248101",
        2764 => x"83244101",
        2765 => x"03290101",
        2766 => x"8329c100",
        2767 => x"032a8100",
        2768 => x"832a4100",
        2769 => x"032b0100",
        2770 => x"13010102",
        2771 => x"67800000",
        2772 => x"13860400",
        2773 => x"13050a00",
        2774 => x"ef001062",
        2775 => x"13090500",
        2776 => x"e31c05f6",
        2777 => x"83250401",
        2778 => x"13050a00",
        2779 => x"eff05fb6",
        2780 => x"9307c000",
        2781 => x"2320fa00",
        2782 => x"8357c400",
        2783 => x"1305f0ff",
        2784 => x"93e70704",
        2785 => x"2316f400",
        2786 => x"6ff01ffa",
        2787 => x"83278600",
        2788 => x"130101fd",
        2789 => x"232e3101",
        2790 => x"23267101",
        2791 => x"23261102",
        2792 => x"23248102",
        2793 => x"23229102",
        2794 => x"23202103",
        2795 => x"232c4101",
        2796 => x"232a5101",
        2797 => x"23286101",
        2798 => x"23248101",
        2799 => x"23229101",
        2800 => x"2320a101",
        2801 => x"832b0600",
        2802 => x"93090600",
        2803 => x"63980712",
        2804 => x"13050000",
        2805 => x"8320c102",
        2806 => x"03248102",
        2807 => x"23a20900",
        2808 => x"83244102",
        2809 => x"03290102",
        2810 => x"8329c101",
        2811 => x"032a8101",
        2812 => x"832a4101",
        2813 => x"032b0101",
        2814 => x"832bc100",
        2815 => x"032c8100",
        2816 => x"832c4100",
        2817 => x"032d0100",
        2818 => x"13010103",
        2819 => x"67800000",
        2820 => x"03ab0b00",
        2821 => x"03ad4b00",
        2822 => x"938b8b00",
        2823 => x"03298400",
        2824 => x"832a0400",
        2825 => x"e3060dfe",
        2826 => x"63642d09",
        2827 => x"8317c400",
        2828 => x"13f70748",
        2829 => x"63020708",
        2830 => x"83244401",
        2831 => x"83250401",
        2832 => x"b3049c02",
        2833 => x"b38aba40",
        2834 => x"13871a00",
        2835 => x"3307a701",
        2836 => x"b3c49403",
        2837 => x"63f4e400",
        2838 => x"93040700",
        2839 => x"93f70740",
        2840 => x"638c070a",
        2841 => x"93850400",
        2842 => x"13050a00",
        2843 => x"eff09fbe",
        2844 => x"13090500",
        2845 => x"6302050c",
        2846 => x"83250401",
        2847 => x"13860a00",
        2848 => x"efd09fa9",
        2849 => x"8357c400",
        2850 => x"93f7f7b7",
        2851 => x"93e70708",
        2852 => x"2316f400",
        2853 => x"23282401",
        2854 => x"232a9400",
        2855 => x"33095901",
        2856 => x"b3845441",
        2857 => x"23202401",
        2858 => x"23249400",
        2859 => x"13090d00",
        2860 => x"63742d01",
        2861 => x"13090d00",
        2862 => x"03250400",
        2863 => x"93050b00",
        2864 => x"13060900",
        2865 => x"efd09fa7",
        2866 => x"83278400",
        2867 => x"330bab01",
        2868 => x"b3872741",
        2869 => x"2324f400",
        2870 => x"83270400",
        2871 => x"b3872701",
        2872 => x"2320f400",
        2873 => x"83a78900",
        2874 => x"b387a741",
        2875 => x"23a4f900",
        2876 => x"e38007ee",
        2877 => x"130d0000",
        2878 => x"6ff05ff2",
        2879 => x"130a0500",
        2880 => x"13840500",
        2881 => x"130b0000",
        2882 => x"130d0000",
        2883 => x"130c3000",
        2884 => x"930c2000",
        2885 => x"6ff09ff0",
        2886 => x"13860400",
        2887 => x"13050a00",
        2888 => x"ef009045",
        2889 => x"13090500",
        2890 => x"e31605f6",
        2891 => x"83250401",
        2892 => x"13050a00",
        2893 => x"eff0df99",
        2894 => x"9307c000",
        2895 => x"2320fa00",
        2896 => x"8357c400",
        2897 => x"1305f0ff",
        2898 => x"93e70704",
        2899 => x"2316f400",
        2900 => x"23a40900",
        2901 => x"6ff01fe8",
        2902 => x"83d7c500",
        2903 => x"130101f6",
        2904 => x"232c8108",
        2905 => x"232a9108",
        2906 => x"23282109",
        2907 => x"23244109",
        2908 => x"232e1108",
        2909 => x"23263109",
        2910 => x"23225109",
        2911 => x"23206109",
        2912 => x"232e7107",
        2913 => x"232c8107",
        2914 => x"232a9107",
        2915 => x"93f70708",
        2916 => x"130a0500",
        2917 => x"13890500",
        2918 => x"93040600",
        2919 => x"13840600",
        2920 => x"63840706",
        2921 => x"83a70501",
        2922 => x"63900706",
        2923 => x"93050004",
        2924 => x"eff05faa",
        2925 => x"2320a900",
        2926 => x"2328a900",
        2927 => x"63120504",
        2928 => x"9307c000",
        2929 => x"2320fa00",
        2930 => x"1305f0ff",
        2931 => x"8320c109",
        2932 => x"03248109",
        2933 => x"83244109",
        2934 => x"03290109",
        2935 => x"8329c108",
        2936 => x"032a8108",
        2937 => x"832a4108",
        2938 => x"032b0108",
        2939 => x"832bc107",
        2940 => x"032c8107",
        2941 => x"832c4107",
        2942 => x"1301010a",
        2943 => x"67800000",
        2944 => x"93070004",
        2945 => x"232af900",
        2946 => x"93070002",
        2947 => x"a304f102",
        2948 => x"93070003",
        2949 => x"23220102",
        2950 => x"2305f102",
        2951 => x"23268100",
        2952 => x"930b5002",
        2953 => x"971a0000",
        2954 => x"938acaf5",
        2955 => x"130c1000",
        2956 => x"130ba000",
        2957 => x"13840400",
        2958 => x"83470400",
        2959 => x"63840700",
        2960 => x"6398770d",
        2961 => x"b30c9440",
        2962 => x"63069402",
        2963 => x"93860c00",
        2964 => x"13860400",
        2965 => x"93050900",
        2966 => x"13050a00",
        2967 => x"eff0dfbc",
        2968 => x"9307f0ff",
        2969 => x"6306f524",
        2970 => x"83274102",
        2971 => x"b3879701",
        2972 => x"2322f102",
        2973 => x"83470400",
        2974 => x"638c0722",
        2975 => x"9307f0ff",
        2976 => x"93041400",
        2977 => x"23280100",
        2978 => x"232e0100",
        2979 => x"232af100",
        2980 => x"232c0100",
        2981 => x"a3090104",
        2982 => x"23240106",
        2983 => x"83c50400",
        2984 => x"13065000",
        2985 => x"13850a00",
        2986 => x"ef009022",
        2987 => x"83270101",
        2988 => x"13841400",
        2989 => x"63120506",
        2990 => x"13f70701",
        2991 => x"63060700",
        2992 => x"13070002",
        2993 => x"a309e104",
        2994 => x"13f78700",
        2995 => x"63060700",
        2996 => x"1307b002",
        2997 => x"a309e104",
        2998 => x"83c60400",
        2999 => x"1307a002",
        3000 => x"6388e604",
        3001 => x"8327c101",
        3002 => x"13840400",
        3003 => x"93060000",
        3004 => x"13069000",
        3005 => x"03470400",
        3006 => x"93051400",
        3007 => x"130707fd",
        3008 => x"637ce608",
        3009 => x"63820604",
        3010 => x"232ef100",
        3011 => x"6f00c003",
        3012 => x"13041400",
        3013 => x"6ff05ff2",
        3014 => x"33055541",
        3015 => x"3315ac00",
        3016 => x"b3e7a700",
        3017 => x"2328f100",
        3018 => x"93040400",
        3019 => x"6ff01ff7",
        3020 => x"0327c100",
        3021 => x"93064700",
        3022 => x"03270700",
        3023 => x"2326d100",
        3024 => x"63420704",
        3025 => x"232ee100",
        3026 => x"03470400",
        3027 => x"9307e002",
        3028 => x"6312f708",
        3029 => x"03471400",
        3030 => x"9307a002",
        3031 => x"6318f704",
        3032 => x"8327c100",
        3033 => x"13042400",
        3034 => x"13874700",
        3035 => x"83a70700",
        3036 => x"2326e100",
        3037 => x"63d40700",
        3038 => x"9307f0ff",
        3039 => x"232af100",
        3040 => x"6f004005",
        3041 => x"3307e040",
        3042 => x"93e72700",
        3043 => x"232ee100",
        3044 => x"2328f100",
        3045 => x"6ff05ffb",
        3046 => x"b3876703",
        3047 => x"13840500",
        3048 => x"93061000",
        3049 => x"b387e700",
        3050 => x"6ff0dff4",
        3051 => x"13041400",
        3052 => x"232a0100",
        3053 => x"93060000",
        3054 => x"93070000",
        3055 => x"13069000",
        3056 => x"03470400",
        3057 => x"93051400",
        3058 => x"130707fd",
        3059 => x"637ae608",
        3060 => x"e39606fa",
        3061 => x"83450400",
        3062 => x"13063000",
        3063 => x"17150000",
        3064 => x"1305c5da",
        3065 => x"ef00d00e",
        3066 => x"63040502",
        3067 => x"97170000",
        3068 => x"9387c7d9",
        3069 => x"3305f540",
        3070 => x"83270101",
        3071 => x"13070004",
        3072 => x"3317a700",
        3073 => x"b3e7e700",
        3074 => x"13041400",
        3075 => x"2328f100",
        3076 => x"83450400",
        3077 => x"13066000",
        3078 => x"17150000",
        3079 => x"130545d7",
        3080 => x"93041400",
        3081 => x"2304b102",
        3082 => x"ef00900a",
        3083 => x"630c0508",
        3084 => x"93070000",
        3085 => x"63980704",
        3086 => x"03270101",
        3087 => x"8327c100",
        3088 => x"13770710",
        3089 => x"63080702",
        3090 => x"93874700",
        3091 => x"2326f100",
        3092 => x"83274102",
        3093 => x"b3873701",
        3094 => x"2322f102",
        3095 => x"6ff09fdd",
        3096 => x"b3876703",
        3097 => x"13840500",
        3098 => x"93061000",
        3099 => x"b387e700",
        3100 => x"6ff01ff5",
        3101 => x"93877700",
        3102 => x"93f787ff",
        3103 => x"93878700",
        3104 => x"6ff0dffc",
        3105 => x"1307c100",
        3106 => x"97060000",
        3107 => x"9386069a",
        3108 => x"13060900",
        3109 => x"93050101",
        3110 => x"13050a00",
        3111 => x"97000000",
        3112 => x"e7000000",
        3113 => x"9307f0ff",
        3114 => x"93090500",
        3115 => x"e312f5fa",
        3116 => x"8357c900",
        3117 => x"93f70704",
        3118 => x"e39807d0",
        3119 => x"03254102",
        3120 => x"6ff0dfd0",
        3121 => x"1307c100",
        3122 => x"97060000",
        3123 => x"93860696",
        3124 => x"13060900",
        3125 => x"93050101",
        3126 => x"13050a00",
        3127 => x"ef00801b",
        3128 => x"6ff05ffc",
        3129 => x"130101fd",
        3130 => x"232a5101",
        3131 => x"83a70501",
        3132 => x"930a0700",
        3133 => x"03a78500",
        3134 => x"23248102",
        3135 => x"23202103",
        3136 => x"232e3101",
        3137 => x"232c4101",
        3138 => x"23261102",
        3139 => x"23229102",
        3140 => x"23286101",
        3141 => x"23267101",
        3142 => x"93090500",
        3143 => x"13840500",
        3144 => x"13090600",
        3145 => x"138a0600",
        3146 => x"63d4e700",
        3147 => x"93070700",
        3148 => x"2320f900",
        3149 => x"03473404",
        3150 => x"63060700",
        3151 => x"93871700",
        3152 => x"2320f900",
        3153 => x"83270400",
        3154 => x"93f70702",
        3155 => x"63880700",
        3156 => x"83270900",
        3157 => x"93872700",
        3158 => x"2320f900",
        3159 => x"83240400",
        3160 => x"93f46400",
        3161 => x"639e0400",
        3162 => x"130b9401",
        3163 => x"930bf0ff",
        3164 => x"8327c400",
        3165 => x"03270900",
        3166 => x"b387e740",
        3167 => x"63c2f408",
        3168 => x"83473404",
        3169 => x"b336f000",
        3170 => x"83270400",
        3171 => x"93f70702",
        3172 => x"6390070c",
        3173 => x"13063404",
        3174 => x"93050a00",
        3175 => x"13850900",
        3176 => x"e7800a00",
        3177 => x"9307f0ff",
        3178 => x"6308f506",
        3179 => x"83270400",
        3180 => x"13074000",
        3181 => x"93040000",
        3182 => x"93f76700",
        3183 => x"639ce700",
        3184 => x"8324c400",
        3185 => x"83270900",
        3186 => x"b384f440",
        3187 => x"63d40400",
        3188 => x"93040000",
        3189 => x"83278400",
        3190 => x"03270401",
        3191 => x"6356f700",
        3192 => x"b387e740",
        3193 => x"b384f400",
        3194 => x"13090000",
        3195 => x"1304a401",
        3196 => x"130bf0ff",
        3197 => x"63902409",
        3198 => x"13050000",
        3199 => x"6f000002",
        3200 => x"93061000",
        3201 => x"13060b00",
        3202 => x"93050a00",
        3203 => x"13850900",
        3204 => x"e7800a00",
        3205 => x"631a7503",
        3206 => x"1305f0ff",
        3207 => x"8320c102",
        3208 => x"03248102",
        3209 => x"83244102",
        3210 => x"03290102",
        3211 => x"8329c101",
        3212 => x"032a8101",
        3213 => x"832a4101",
        3214 => x"032b0101",
        3215 => x"832bc100",
        3216 => x"13010103",
        3217 => x"67800000",
        3218 => x"93841400",
        3219 => x"6ff05ff2",
        3220 => x"3307d400",
        3221 => x"13060003",
        3222 => x"a301c704",
        3223 => x"03475404",
        3224 => x"93871600",
        3225 => x"b307f400",
        3226 => x"93862600",
        3227 => x"a381e704",
        3228 => x"6ff05ff2",
        3229 => x"93061000",
        3230 => x"13060400",
        3231 => x"93050a00",
        3232 => x"13850900",
        3233 => x"e7800a00",
        3234 => x"e30865f9",
        3235 => x"13091900",
        3236 => x"6ff05ff6",
        3237 => x"130101fd",
        3238 => x"23248102",
        3239 => x"23229102",
        3240 => x"23202103",
        3241 => x"232e3101",
        3242 => x"23261102",
        3243 => x"232c4101",
        3244 => x"232a5101",
        3245 => x"23286101",
        3246 => x"03c88501",
        3247 => x"93078007",
        3248 => x"93040500",
        3249 => x"13840500",
        3250 => x"13090600",
        3251 => x"93890600",
        3252 => x"63e20703",
        3253 => x"93072006",
        3254 => x"93863504",
        3255 => x"63e20703",
        3256 => x"63040828",
        3257 => x"93078005",
        3258 => x"17160000",
        3259 => x"1306c6aa",
        3260 => x"630cf81c",
        3261 => x"930a2404",
        3262 => x"23010405",
        3263 => x"6f008004",
        3264 => x"9307d8f9",
        3265 => x"93f7f70f",
        3266 => x"13065001",
        3267 => x"e364f6fe",
        3268 => x"17160000",
        3269 => x"1306c6ba",
        3270 => x"93972700",
        3271 => x"b387c700",
        3272 => x"83a70700",
        3273 => x"b387c700",
        3274 => x"67800700",
        3275 => x"83270700",
        3276 => x"938a2504",
        3277 => x"93864700",
        3278 => x"83a70700",
        3279 => x"2320d700",
        3280 => x"2381f504",
        3281 => x"93071000",
        3282 => x"6f00c025",
        3283 => x"83a70500",
        3284 => x"03250700",
        3285 => x"13f60708",
        3286 => x"93054500",
        3287 => x"63060602",
        3288 => x"83270500",
        3289 => x"2320b700",
        3290 => x"63d80700",
        3291 => x"1307d002",
        3292 => x"b307f040",
        3293 => x"a301e404",
        3294 => x"17160000",
        3295 => x"1306c6a1",
        3296 => x"1308a000",
        3297 => x"6f004006",
        3298 => x"13f60704",
        3299 => x"83270500",
        3300 => x"2320b700",
        3301 => x"e30a06fc",
        3302 => x"93970701",
        3303 => x"93d70741",
        3304 => x"6ff09ffc",
        3305 => x"83a50500",
        3306 => x"03260700",
        3307 => x"13f50508",
        3308 => x"83270600",
        3309 => x"13064600",
        3310 => x"631a0500",
        3311 => x"93f50504",
        3312 => x"63860500",
        3313 => x"93970701",
        3314 => x"93d70701",
        3315 => x"2320c700",
        3316 => x"1307f006",
        3317 => x"17160000",
        3318 => x"1306069c",
        3319 => x"6314e814",
        3320 => x"13088000",
        3321 => x"a3010404",
        3322 => x"03274400",
        3323 => x"2324e400",
        3324 => x"634e0700",
        3325 => x"83250400",
        3326 => x"33e7e700",
        3327 => x"938a0600",
        3328 => x"93f5b5ff",
        3329 => x"2320b400",
        3330 => x"63040702",
        3331 => x"938a0600",
        3332 => x"33f70703",
        3333 => x"938afaff",
        3334 => x"3307e600",
        3335 => x"03470700",
        3336 => x"2380ea00",
        3337 => x"13870700",
        3338 => x"b3d70703",
        3339 => x"e37207ff",
        3340 => x"93078000",
        3341 => x"6314f802",
        3342 => x"83270400",
        3343 => x"93f71700",
        3344 => x"638e0700",
        3345 => x"03274400",
        3346 => x"83270401",
        3347 => x"63c8e700",
        3348 => x"93070003",
        3349 => x"a38ffafe",
        3350 => x"938afaff",
        3351 => x"b3865641",
        3352 => x"2328d400",
        3353 => x"13870900",
        3354 => x"93060900",
        3355 => x"1306c100",
        3356 => x"93050400",
        3357 => x"13850400",
        3358 => x"eff0dfc6",
        3359 => x"130af0ff",
        3360 => x"63184513",
        3361 => x"1305f0ff",
        3362 => x"8320c102",
        3363 => x"03248102",
        3364 => x"83244102",
        3365 => x"03290102",
        3366 => x"8329c101",
        3367 => x"032a8101",
        3368 => x"832a4101",
        3369 => x"032b0101",
        3370 => x"13010103",
        3371 => x"67800000",
        3372 => x"83a70500",
        3373 => x"93e70702",
        3374 => x"23a0f500",
        3375 => x"13088007",
        3376 => x"17160000",
        3377 => x"1306868e",
        3378 => x"a3020405",
        3379 => x"83250400",
        3380 => x"03250700",
        3381 => x"13f80508",
        3382 => x"83270500",
        3383 => x"13054500",
        3384 => x"631a0800",
        3385 => x"13f80504",
        3386 => x"63060800",
        3387 => x"93970701",
        3388 => x"93d70701",
        3389 => x"2320a700",
        3390 => x"13f71500",
        3391 => x"63060700",
        3392 => x"93e50502",
        3393 => x"2320b400",
        3394 => x"63860700",
        3395 => x"13080001",
        3396 => x"6ff05fed",
        3397 => x"03270400",
        3398 => x"1377f7fd",
        3399 => x"2320e400",
        3400 => x"6ff0dffe",
        3401 => x"1308a000",
        3402 => x"6ff0dfeb",
        3403 => x"03a60500",
        3404 => x"83270700",
        3405 => x"83a54501",
        3406 => x"13780608",
        3407 => x"13854700",
        3408 => x"630a0800",
        3409 => x"2320a700",
        3410 => x"83a70700",
        3411 => x"23a0b700",
        3412 => x"6f008001",
        3413 => x"2320a700",
        3414 => x"13760604",
        3415 => x"83a70700",
        3416 => x"e30606fe",
        3417 => x"2390b700",
        3418 => x"23280400",
        3419 => x"938a0600",
        3420 => x"6ff05fef",
        3421 => x"83270700",
        3422 => x"03a64500",
        3423 => x"93050000",
        3424 => x"93864700",
        3425 => x"2320d700",
        3426 => x"83aa0700",
        3427 => x"13850a00",
        3428 => x"ef000034",
        3429 => x"63060500",
        3430 => x"33055541",
        3431 => x"2322a400",
        3432 => x"83274400",
        3433 => x"2328f400",
        3434 => x"a3010404",
        3435 => x"6ff09feb",
        3436 => x"83260401",
        3437 => x"13860a00",
        3438 => x"93050900",
        3439 => x"13850400",
        3440 => x"e7800900",
        3441 => x"e30045ed",
        3442 => x"83270400",
        3443 => x"93f72700",
        3444 => x"63940704",
        3445 => x"8327c100",
        3446 => x"0325c400",
        3447 => x"e356f5ea",
        3448 => x"13850700",
        3449 => x"6ff05fea",
        3450 => x"93061000",
        3451 => x"13860a00",
        3452 => x"93050900",
        3453 => x"13850400",
        3454 => x"e7800900",
        3455 => x"e30465e9",
        3456 => x"130a1a00",
        3457 => x"8327c400",
        3458 => x"0327c100",
        3459 => x"b387e740",
        3460 => x"e34cfafc",
        3461 => x"6ff01ffc",
        3462 => x"130a0000",
        3463 => x"930a9401",
        3464 => x"130bf0ff",
        3465 => x"6ff01ffe",
        3466 => x"8397c500",
        3467 => x"130101fe",
        3468 => x"232c8100",
        3469 => x"232a9100",
        3470 => x"232e1100",
        3471 => x"23282101",
        3472 => x"23263101",
        3473 => x"13f78700",
        3474 => x"93040500",
        3475 => x"13840500",
        3476 => x"631a0712",
        3477 => x"03a74500",
        3478 => x"6346e000",
        3479 => x"03a70504",
        3480 => x"6356e010",
        3481 => x"0327c402",
        3482 => x"63020710",
        3483 => x"03a90400",
        3484 => x"93963701",
        3485 => x"23a00400",
        3486 => x"83250402",
        3487 => x"63dc060a",
        3488 => x"03264405",
        3489 => x"8357c400",
        3490 => x"93f74700",
        3491 => x"638e0700",
        3492 => x"83274400",
        3493 => x"3306f640",
        3494 => x"83274403",
        3495 => x"63860700",
        3496 => x"83270404",
        3497 => x"3306f640",
        3498 => x"8327c402",
        3499 => x"83250402",
        3500 => x"93060000",
        3501 => x"13850400",
        3502 => x"e7800700",
        3503 => x"1307f0ff",
        3504 => x"8357c400",
        3505 => x"6312e502",
        3506 => x"83a60400",
        3507 => x"1307d001",
        3508 => x"6362d70a",
        3509 => x"37074020",
        3510 => x"13071700",
        3511 => x"3357d700",
        3512 => x"13771700",
        3513 => x"63080708",
        3514 => x"03270401",
        3515 => x"23220400",
        3516 => x"2320e400",
        3517 => x"13973701",
        3518 => x"635c0700",
        3519 => x"9307f0ff",
        3520 => x"6316f500",
        3521 => x"83a70400",
        3522 => x"63940700",
        3523 => x"232aa404",
        3524 => x"83254403",
        3525 => x"23a02401",
        3526 => x"638a0504",
        3527 => x"93074404",
        3528 => x"6386f500",
        3529 => x"13850400",
        3530 => x"efe09ffa",
        3531 => x"232a0402",
        3532 => x"6f00c003",
        3533 => x"13060000",
        3534 => x"93061000",
        3535 => x"13850400",
        3536 => x"e7000700",
        3537 => x"9307f0ff",
        3538 => x"13060500",
        3539 => x"e31cf5f2",
        3540 => x"83a70400",
        3541 => x"e38807f2",
        3542 => x"1307d001",
        3543 => x"6386e700",
        3544 => x"13076001",
        3545 => x"6394e706",
        3546 => x"23a02401",
        3547 => x"13050000",
        3548 => x"6f00c006",
        3549 => x"93e70704",
        3550 => x"93970701",
        3551 => x"93d70741",
        3552 => x"6f004005",
        3553 => x"83a90501",
        3554 => x"e38209fe",
        3555 => x"03a90500",
        3556 => x"93f73700",
        3557 => x"23a03501",
        3558 => x"33093941",
        3559 => x"13070000",
        3560 => x"63940700",
        3561 => x"03a74501",
        3562 => x"2324e400",
        3563 => x"e35020fd",
        3564 => x"83278402",
        3565 => x"83250402",
        3566 => x"93060900",
        3567 => x"13860900",
        3568 => x"13850400",
        3569 => x"e7800700",
        3570 => x"6348a002",
        3571 => x"8317c400",
        3572 => x"93e70704",
        3573 => x"2316f400",
        3574 => x"1305f0ff",
        3575 => x"8320c101",
        3576 => x"03248101",
        3577 => x"83244101",
        3578 => x"03290101",
        3579 => x"8329c100",
        3580 => x"13010102",
        3581 => x"67800000",
        3582 => x"b389a900",
        3583 => x"3309a940",
        3584 => x"6ff0dffa",
        3585 => x"83a70501",
        3586 => x"130101ff",
        3587 => x"23261100",
        3588 => x"23248100",
        3589 => x"23229100",
        3590 => x"63900702",
        3591 => x"93040000",
        3592 => x"8320c100",
        3593 => x"03248100",
        3594 => x"13850400",
        3595 => x"83244100",
        3596 => x"13010101",
        3597 => x"67800000",
        3598 => x"93040500",
        3599 => x"13840500",
        3600 => x"63080500",
        3601 => x"83270502",
        3602 => x"63940700",
        3603 => x"efe00ffe",
        3604 => x"8317c400",
        3605 => x"e38407fc",
        3606 => x"03274406",
        3607 => x"13771700",
        3608 => x"631a0700",
        3609 => x"93f70720",
        3610 => x"63960700",
        3611 => x"03258405",
        3612 => x"efe05fe3",
        3613 => x"13850400",
        3614 => x"93050400",
        3615 => x"eff0dfda",
        3616 => x"83274406",
        3617 => x"93040500",
        3618 => x"93f71700",
        3619 => x"e39a07f8",
        3620 => x"8357c400",
        3621 => x"93f70720",
        3622 => x"e39407f8",
        3623 => x"03258405",
        3624 => x"efe0dfe1",
        3625 => x"6ff0dff7",
        3626 => x"93050500",
        3627 => x"631e0500",
        3628 => x"13868181",
        3629 => x"97050000",
        3630 => x"938505f5",
        3631 => x"17c5ff1f",
        3632 => x"13058576",
        3633 => x"6fe01f80",
        3634 => x"03a54187",
        3635 => x"6ff09ff3",
        3636 => x"93f5f50f",
        3637 => x"3306c500",
        3638 => x"6316c500",
        3639 => x"13050000",
        3640 => x"67800000",
        3641 => x"83470500",
        3642 => x"e38cb7fe",
        3643 => x"13051500",
        3644 => x"6ff09ffe",
        3645 => x"130101ff",
        3646 => x"23248100",
        3647 => x"13040500",
        3648 => x"13850500",
        3649 => x"93050600",
        3650 => x"23a20188",
        3651 => x"23261100",
        3652 => x"efc0dfe6",
        3653 => x"9307f0ff",
        3654 => x"6318f500",
        3655 => x"83a74188",
        3656 => x"63840700",
        3657 => x"2320f400",
        3658 => x"8320c100",
        3659 => x"03248100",
        3660 => x"13010101",
        3661 => x"67800000",
        3662 => x"130101ff",
        3663 => x"23248100",
        3664 => x"13040500",
        3665 => x"13850500",
        3666 => x"23a20188",
        3667 => x"23261100",
        3668 => x"efd08f8a",
        3669 => x"9307f0ff",
        3670 => x"6318f500",
        3671 => x"83a74188",
        3672 => x"63840700",
        3673 => x"2320f400",
        3674 => x"8320c100",
        3675 => x"03248100",
        3676 => x"13010101",
        3677 => x"67800000",
        3678 => x"130101fe",
        3679 => x"232c8100",
        3680 => x"232e1100",
        3681 => x"232a9100",
        3682 => x"23282101",
        3683 => x"23263101",
        3684 => x"23244101",
        3685 => x"13040600",
        3686 => x"63940502",
        3687 => x"03248101",
        3688 => x"8320c101",
        3689 => x"83244101",
        3690 => x"03290101",
        3691 => x"8329c100",
        3692 => x"032a8100",
        3693 => x"93050600",
        3694 => x"13010102",
        3695 => x"6fe09fe9",
        3696 => x"63180602",
        3697 => x"efe0dfd0",
        3698 => x"93040000",
        3699 => x"8320c101",
        3700 => x"03248101",
        3701 => x"03290101",
        3702 => x"8329c100",
        3703 => x"032a8100",
        3704 => x"13850400",
        3705 => x"83244101",
        3706 => x"13010102",
        3707 => x"67800000",
        3708 => x"130a0500",
        3709 => x"93840500",
        3710 => x"ef008005",
        3711 => x"13090500",
        3712 => x"63668500",
        3713 => x"93571500",
        3714 => x"e3e287fc",
        3715 => x"93050400",
        3716 => x"13050a00",
        3717 => x"efe01fe4",
        3718 => x"93090500",
        3719 => x"63160500",
        3720 => x"93840900",
        3721 => x"6ff09ffa",
        3722 => x"13060400",
        3723 => x"63748900",
        3724 => x"13060900",
        3725 => x"93850400",
        3726 => x"13850900",
        3727 => x"efc0dfcd",
        3728 => x"93850400",
        3729 => x"13050a00",
        3730 => x"efe09fc8",
        3731 => x"6ff05ffd",
        3732 => x"83a7c5ff",
        3733 => x"1385c7ff",
        3734 => x"63d80700",
        3735 => x"b385a500",
        3736 => x"83a70500",
        3737 => x"3305f500",
        3738 => x"67800000",
        3739 => x"10000000",
        3740 => x"00000000",
        3741 => x"037a5200",
        3742 => x"017c0101",
        3743 => x"1b0d0200",
        3744 => x"10000000",
        3745 => x"18000000",
        3746 => x"20d4ffff",
        3747 => x"fc040000",
        3748 => x"00000000",
        3749 => x"10000000",
        3750 => x"00000000",
        3751 => x"037a5200",
        3752 => x"017c0101",
        3753 => x"1b0d0200",
        3754 => x"10000000",
        3755 => x"18000000",
        3756 => x"f4d8ffff",
        3757 => x"b0040000",
        3758 => x"00000000",
        3759 => x"10000000",
        3760 => x"00000000",
        3761 => x"037a5200",
        3762 => x"017c0101",
        3763 => x"1b0d0200",
        3764 => x"10000000",
        3765 => x"18000000",
        3766 => x"7cddffff",
        3767 => x"70040000",
        3768 => x"00000000",
        3769 => x"30313233",
        3770 => x"34353637",
        3771 => x"38396162",
        3772 => x"63646566",
        3773 => x"00000000",
        3774 => x"a4040000",
        3775 => x"dc030000",
        3776 => x"dc030000",
        3777 => x"dc030000",
        3778 => x"b0040000",
        3779 => x"dc030000",
        3780 => x"dc030000",
        3781 => x"dc030000",
        3782 => x"dc030000",
        3783 => x"dc030000",
        3784 => x"dc030000",
        3785 => x"dc030000",
        3786 => x"dc030000",
        3787 => x"dc030000",
        3788 => x"dc030000",
        3789 => x"bc040000",
        3790 => x"dc030000",
        3791 => x"c8040000",
        3792 => x"d4040000",
        3793 => x"dc030000",
        3794 => x"e0040000",
        3795 => x"ec040000",
        3796 => x"dc030000",
        3797 => x"f8040000",
        3798 => x"98040000",
        3799 => x"dc030000",
        3800 => x"dc030000",
        3801 => x"dc030000",
        3802 => x"04050000",
        3803 => x"dc030000",
        3804 => x"dc030000",
        3805 => x"dc030000",
        3806 => x"dc030000",
        3807 => x"dc030000",
        3808 => x"dc030000",
        3809 => x"dc030000",
        3810 => x"14050000",
        3811 => x"a8050000",
        3812 => x"c0050000",
        3813 => x"f0050000",
        3814 => x"70050000",
        3815 => x"70050000",
        3816 => x"70050000",
        3817 => x"70050000",
        3818 => x"70050000",
        3819 => x"70050000",
        3820 => x"d8050000",
        3821 => x"70050000",
        3822 => x"70050000",
        3823 => x"70050000",
        3824 => x"70050000",
        3825 => x"88050000",
        3826 => x"88050000",
        3827 => x"a8050000",
        3828 => x"70050000",
        3829 => x"70050000",
        3830 => x"70050000",
        3831 => x"70050000",
        3832 => x"9c050000",
        3833 => x"08060000",
        3834 => x"30060000",
        3835 => x"70050000",
        3836 => x"70050000",
        3837 => x"70050000",
        3838 => x"70050000",
        3839 => x"70050000",
        3840 => x"70050000",
        3841 => x"70050000",
        3842 => x"70050000",
        3843 => x"70050000",
        3844 => x"70050000",
        3845 => x"70050000",
        3846 => x"70050000",
        3847 => x"70050000",
        3848 => x"70050000",
        3849 => x"88050000",
        3850 => x"88050000",
        3851 => x"70050000",
        3852 => x"70050000",
        3853 => x"70050000",
        3854 => x"70050000",
        3855 => x"70050000",
        3856 => x"70050000",
        3857 => x"70050000",
        3858 => x"70050000",
        3859 => x"70050000",
        3860 => x"70050000",
        3861 => x"70050000",
        3862 => x"70050000",
        3863 => x"9c050000",
        3864 => x"0d0a4542",
        3865 => x"5245414b",
        3866 => x"21206d65",
        3867 => x"7063203d",
        3868 => x"20000000",
        3869 => x"20696e73",
        3870 => x"6e203d20",
        3871 => x"00000000",
        3872 => x"0d0a0000",
        3873 => x"0d0a0a44",
        3874 => x"6973706c",
        3875 => x"6179696e",
        3876 => x"67207468",
        3877 => x"65207469",
        3878 => x"6d652070",
        3879 => x"61737365",
        3880 => x"64207369",
        3881 => x"6e636520",
        3882 => x"72657365",
        3883 => x"740d0a0a",
        3884 => x"00000000",
        3885 => x"2530356c",
        3886 => x"643a2530",
        3887 => x"366c6420",
        3888 => x"20202530",
        3889 => x"326c643a",
        3890 => x"2530326c",
        3891 => x"643a2530",
        3892 => x"326c640d",
        3893 => x"00000000",
        3894 => x"696e7465",
        3895 => x"72727570",
        3896 => x"745f6469",
        3897 => x"72656374",
        3898 => x"00000000",
        3899 => x"54485541",
        3900 => x"53205249",
        3901 => x"53432d56",
        3902 => x"20525633",
        3903 => x"32494d20",
        3904 => x"62617265",
        3905 => x"206d6574",
        3906 => x"616c2070",
        3907 => x"726f6365",
        3908 => x"73736f72",
        3909 => x"00000000",
        3910 => x"54686520",
        3911 => x"48616775",
        3912 => x"6520556e",
        3913 => x"69766572",
        3914 => x"73697479",
        3915 => x"206f6620",
        3916 => x"4170706c",
        3917 => x"69656420",
        3918 => x"53636965",
        3919 => x"6e636573",
        3920 => x"00000000",
        3921 => x"44657061",
        3922 => x"72746d65",
        3923 => x"6e74206f",
        3924 => x"6620456c",
        3925 => x"65637472",
        3926 => x"6963616c",
        3927 => x"20456e67",
        3928 => x"696e6565",
        3929 => x"72696e67",
        3930 => x"00000000",
        3931 => x"4a2e452e",
        3932 => x"4a2e206f",
        3933 => x"70206465",
        3934 => x"6e204272",
        3935 => x"6f757700",
        3936 => x"232d302b",
        3937 => x"20000000",
        3938 => x"686c4c00",
        3939 => x"65666745",
        3940 => x"46470000",
        3941 => x"30313233",
        3942 => x"34353637",
        3943 => x"38394142",
        3944 => x"43444546",
        3945 => x"00000000",
        3946 => x"30313233",
        3947 => x"34353637",
        3948 => x"38396162",
        3949 => x"63646566",
        3950 => x"00000000",
        3951 => x"00010202",
        3952 => x"03030303",
        3953 => x"04040404",
        3954 => x"04040404",
        3955 => x"05050505",
        3956 => x"05050505",
        3957 => x"05050505",
        3958 => x"05050505",
        3959 => x"06060606",
        3960 => x"06060606",
        3961 => x"06060606",
        3962 => x"06060606",
        3963 => x"06060606",
        3964 => x"06060606",
        3965 => x"06060606",
        3966 => x"06060606",
        3967 => x"07070707",
        3968 => x"07070707",
        3969 => x"07070707",
        3970 => x"07070707",
        3971 => x"07070707",
        3972 => x"07070707",
        3973 => x"07070707",
        3974 => x"07070707",
        3975 => x"07070707",
        3976 => x"07070707",
        3977 => x"07070707",
        3978 => x"07070707",
        3979 => x"07070707",
        3980 => x"07070707",
        3981 => x"07070707",
        3982 => x"07070707",
        3983 => x"08080808",
        3984 => x"08080808",
        3985 => x"08080808",
        3986 => x"08080808",
        3987 => x"08080808",
        3988 => x"08080808",
        3989 => x"08080808",
        3990 => x"08080808",
        3991 => x"08080808",
        3992 => x"08080808",
        3993 => x"08080808",
        3994 => x"08080808",
        3995 => x"08080808",
        3996 => x"08080808",
        3997 => x"08080808",
        3998 => x"08080808",
        3999 => x"08080808",
        4000 => x"08080808",
        4001 => x"08080808",
        4002 => x"08080808",
        4003 => x"08080808",
        4004 => x"08080808",
        4005 => x"08080808",
        4006 => x"08080808",
        4007 => x"08080808",
        4008 => x"08080808",
        4009 => x"08080808",
        4010 => x"08080808",
        4011 => x"08080808",
        4012 => x"08080808",
        4013 => x"08080808",
        4014 => x"08080808",
        4015 => x"70f4ffff",
        4016 => x"90f4ffff",
        4017 => x"38f4ffff",
        4018 => x"38f4ffff",
        4019 => x"38f4ffff",
        4020 => x"38f4ffff",
        4021 => x"90f4ffff",
        4022 => x"38f4ffff",
        4023 => x"38f4ffff",
        4024 => x"38f4ffff",
        4025 => x"38f4ffff",
        4026 => x"70f6ffff",
        4027 => x"e8f4ffff",
        4028 => x"f4f5ffff",
        4029 => x"38f4ffff",
        4030 => x"38f4ffff",
        4031 => x"b8f6ffff",
        4032 => x"38f4ffff",
        4033 => x"e8f4ffff",
        4034 => x"38f4ffff",
        4035 => x"38f4ffff",
        4036 => x"00f6ffff",
        4037 => x"d83c0000",
        4038 => x"ec3c0000",
        4039 => x"183d0000",
        4040 => x"443d0000",
        4041 => x"6c3d0000",
        4042 => x"00000000",
        4043 => x"00000000",
        4044 => x"03000000",
        4045 => x"b0000020",
        4046 => x"00000000",
        4047 => x"b0000020",
        4048 => x"18010020",
        4049 => x"80010020",
        4050 => x"00000000",
        4051 => x"00000000",
        4052 => x"00000000",
        4053 => x"00000000",
        4054 => x"00000000",
        4055 => x"00000000",
        4056 => x"00000000",
        4057 => x"00000000",
        4058 => x"00000000",
        4059 => x"00000000",
        4060 => x"00000000",
        4061 => x"00000000",
        4062 => x"00000000",
        4063 => x"00000000",
        4064 => x"00000000",
        4065 => x"78000020",
        4066 => x"24000020",
        4067 => x"00000000"
            );
end package rom_image;
