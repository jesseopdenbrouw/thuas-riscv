-- srec2vhdl table generator
-- for input file 'bootloader.srec'
-- date: Mon Jan 15 17:30:46 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package bootrom_image is
    constant bootrom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382c255",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"b7070020",
           9 => x"93870700",
          10 => x"13070500",
          11 => x"3386e740",
          12 => x"63f4e700",
          13 => x"13060000",
          14 => x"93050000",
          15 => x"13050500",
          16 => x"ef000052",
          17 => x"37050020",
          18 => x"b7070020",
          19 => x"93870700",
          20 => x"13070500",
          21 => x"3386e740",
          22 => x"63f4e700",
          23 => x"13060000",
          24 => x"b7150010",
          25 => x"9385c5e1",
          26 => x"13050500",
          27 => x"ef000051",
          28 => x"ef005021",
          29 => x"37c50100",
          30 => x"93050000",
          31 => x"13050520",
          32 => x"ef000070",
          33 => x"37150010",
          34 => x"130585cb",
          35 => x"ef000074",
          36 => x"37150010",
          37 => x"1305c5cd",
          38 => x"ef004073",
          39 => x"732510fc",
          40 => x"37190010",
          41 => x"ef00500e",
          42 => x"130589cd",
          43 => x"ef000072",
          44 => x"b70700f0",
          45 => x"1307f03f",
          46 => x"370a1000",
          47 => x"b709a000",
          48 => x"23a2e700",
          49 => x"93041000",
          50 => x"130afaff",
          51 => x"b70a00f0",
          52 => x"93891900",
          53 => x"b3f74401",
          54 => x"639c0700",
          55 => x"1305a002",
          56 => x"ef00c06c",
          57 => x"83a74a00",
          58 => x"93d71700",
          59 => x"23a2fa00",
          60 => x"ef00004d",
          61 => x"13040500",
          62 => x"63160504",
          63 => x"93841400",
          64 => x"e39a34fd",
          65 => x"b70700f0",
          66 => x"23a20700",
          67 => x"631a0400",
          68 => x"93050000",
          69 => x"13050000",
          70 => x"ef008066",
          71 => x"e7000400",
          72 => x"ef00004b",
          73 => x"1375f50f",
          74 => x"93071002",
          75 => x"6300f502",
          76 => x"93074002",
          77 => x"93040000",
          78 => x"6316f520",
          79 => x"13041000",
          80 => x"6f00c001",
          81 => x"13041000",
          82 => x"6ff0dffb",
          83 => x"37150010",
          84 => x"130505cf",
          85 => x"ef008067",
          86 => x"13040000",
          87 => x"93040000",
          88 => x"370a00f0",
          89 => x"130b3005",
          90 => x"930ba004",
          91 => x"130c3002",
          92 => x"93092000",
          93 => x"930ca000",
          94 => x"b71a0010",
          95 => x"83274a00",
          96 => x"93c71700",
          97 => x"2322fa00",
          98 => x"ef008044",
          99 => x"1375f50f",
         100 => x"631e6517",
         101 => x"ef00c043",
         102 => x"137df50f",
         103 => x"9307fdfc",
         104 => x"93f7f70f",
         105 => x"63e6f910",
         106 => x"93071003",
         107 => x"631afd04",
         108 => x"13052000",
         109 => x"ef008065",
         110 => x"930dd5ff",
         111 => x"13054000",
         112 => x"ef00c064",
         113 => x"b70601ff",
         114 => x"b705ffff",
         115 => x"130d0500",
         116 => x"b38dad00",
         117 => x"9386f6ff",
         118 => x"9385f50f",
         119 => x"6398ad05",
         120 => x"130da000",
         121 => x"ef00c03e",
         122 => x"1375f50f",
         123 => x"e31ca5ff",
         124 => x"e31604f8",
         125 => x"13850acf",
         126 => x"ef00405d",
         127 => x"6ff01ff8",
         128 => x"93072003",
         129 => x"13052000",
         130 => x"631afd00",
         131 => x"ef000060",
         132 => x"930dc5ff",
         133 => x"13056000",
         134 => x"6ff09ffa",
         135 => x"ef00005f",
         136 => x"930db5ff",
         137 => x"13058000",
         138 => x"6ff09ff9",
         139 => x"1378cdff",
         140 => x"13052000",
         141 => x"2326b100",
         142 => x"2324d100",
         143 => x"23220101",
         144 => x"ef00c05c",
         145 => x"03284100",
         146 => x"93070500",
         147 => x"37060001",
         148 => x"13753d00",
         149 => x"03270800",
         150 => x"83268100",
         151 => x"8325c100",
         152 => x"93083000",
         153 => x"1306f6ff",
         154 => x"13031000",
         155 => x"63063503",
         156 => x"630a1503",
         157 => x"630c6500",
         158 => x"137707f0",
         159 => x"b3e7e700",
         160 => x"2320f800",
         161 => x"130d1d00",
         162 => x"6ff05ff5",
         163 => x"3377b700",
         164 => x"93978700",
         165 => x"6ff09ffe",
         166 => x"3377d700",
         167 => x"93970701",
         168 => x"6ff0dffd",
         169 => x"3377c700",
         170 => x"93978701",
         171 => x"6ff01ffd",
         172 => x"93079dfc",
         173 => x"93f7f70f",
         174 => x"63e2f904",
         175 => x"13052000",
         176 => x"ef00c054",
         177 => x"93077003",
         178 => x"13058000",
         179 => x"630afd00",
         180 => x"93078003",
         181 => x"13056000",
         182 => x"6304fd00",
         183 => x"13054000",
         184 => x"ef00c052",
         185 => x"93040500",
         186 => x"130da000",
         187 => x"ef00402e",
         188 => x"1375f50f",
         189 => x"e31ca5ff",
         190 => x"6ff09fef",
         191 => x"ef00402d",
         192 => x"1375f50f",
         193 => x"e31c95ff",
         194 => x"6ff09fee",
         195 => x"63187509",
         196 => x"63180400",
         197 => x"37150010",
         198 => x"130505cf",
         199 => x"ef00004b",
         200 => x"93050000",
         201 => x"13050000",
         202 => x"ef008045",
         203 => x"b70700f0",
         204 => x"23a20700",
         205 => x"e7800400",
         206 => x"b70700f0",
         207 => x"1307a00a",
         208 => x"23a2e700",
         209 => x"130589cd",
         210 => x"b7190010",
         211 => x"ef000048",
         212 => x"13040000",
         213 => x"b71b0010",
         214 => x"938999ba",
         215 => x"b7170010",
         216 => x"138547cf",
         217 => x"ef008046",
         218 => x"93059002",
         219 => x"13054101",
         220 => x"ef000028",
         221 => x"b7170010",
         222 => x"130a0500",
         223 => x"938587cf",
         224 => x"13054101",
         225 => x"ef00c021",
         226 => x"631e0500",
         227 => x"37150010",
         228 => x"1305c5cf",
         229 => x"ef008043",
         230 => x"6f004003",
         231 => x"e31a85e5",
         232 => x"6ff09ff9",
         233 => x"b7170010",
         234 => x"938587de",
         235 => x"13054101",
         236 => x"ef00001f",
         237 => x"63100502",
         238 => x"93050000",
         239 => x"ef00403c",
         240 => x"b70700f0",
         241 => x"23a20700",
         242 => x"e7800400",
         243 => x"e3080af8",
         244 => x"6f000018",
         245 => x"b7170010",
         246 => x"13063000",
         247 => x"9385c7de",
         248 => x"13054101",
         249 => x"ef00c073",
         250 => x"63100504",
         251 => x"93050000",
         252 => x"13057101",
         253 => x"ef00c04d",
         254 => x"93773500",
         255 => x"13040500",
         256 => x"63960706",
         257 => x"93058000",
         258 => x"ef000061",
         259 => x"37150010",
         260 => x"130505df",
         261 => x"ef00803b",
         262 => x"03250400",
         263 => x"93058000",
         264 => x"ef00805f",
         265 => x"6ff09ffa",
         266 => x"b7170010",
         267 => x"13063000",
         268 => x"9385c7e0",
         269 => x"13054101",
         270 => x"ef00806e",
         271 => x"631e0502",
         272 => x"93050101",
         273 => x"13057101",
         274 => x"ef008048",
         275 => x"93773500",
         276 => x"13040500",
         277 => x"639c0700",
         278 => x"03250101",
         279 => x"93050000",
         280 => x"ef000047",
         281 => x"2320a400",
         282 => x"6ff05ff6",
         283 => x"37150010",
         284 => x"130545df",
         285 => x"6ff01ff2",
         286 => x"13063000",
         287 => x"93850be1",
         288 => x"13054101",
         289 => x"ef00c069",
         290 => x"83474101",
         291 => x"1307e006",
         292 => x"63080508",
         293 => x"6396e70a",
         294 => x"93773400",
         295 => x"e39807fc",
         296 => x"130c0404",
         297 => x"b71c0010",
         298 => x"371d0010",
         299 => x"930d80ff",
         300 => x"93058000",
         301 => x"13050400",
         302 => x"ef000056",
         303 => x"13850cdf",
         304 => x"ef00c030",
         305 => x"032a0400",
         306 => x"93058000",
         307 => x"930a8001",
         308 => x"13050a00",
         309 => x"ef004054",
         310 => x"13054de1",
         311 => x"ef00002f",
         312 => x"370b00ff",
         313 => x"33756a01",
         314 => x"33555501",
         315 => x"b3063501",
         316 => x"83c60600",
         317 => x"93f67609",
         318 => x"63800604",
         319 => x"938a8aff",
         320 => x"ef00c02a",
         321 => x"135b8b00",
         322 => x"e39ebafd",
         323 => x"13044400",
         324 => x"130589cd",
         325 => x"ef00802b",
         326 => x"e31c8cf8",
         327 => x"6ff01fe4",
         328 => x"e38ce7f6",
         329 => x"93050000",
         330 => x"13057101",
         331 => x"ef00403a",
         332 => x"13040500",
         333 => x"6ff05ff6",
         334 => x"1305e002",
         335 => x"6ff01ffc",
         336 => x"e30e0ae0",
         337 => x"37150010",
         338 => x"130585e1",
         339 => x"ef000028",
         340 => x"130589cd",
         341 => x"ef008027",
         342 => x"6ff05fe0",
         343 => x"6f000000",
         344 => x"13030500",
         345 => x"630a0600",
         346 => x"2300b300",
         347 => x"1306f6ff",
         348 => x"13031300",
         349 => x"e31a06fe",
         350 => x"67800000",
         351 => x"13030500",
         352 => x"630e0600",
         353 => x"83830500",
         354 => x"23007300",
         355 => x"1306f6ff",
         356 => x"13031300",
         357 => x"93851500",
         358 => x"e31606fe",
         359 => x"67800000",
         360 => x"03460500",
         361 => x"83c60500",
         362 => x"13051500",
         363 => x"93851500",
         364 => x"6314d600",
         365 => x"e31606fe",
         366 => x"3305d640",
         367 => x"67800000",
         368 => x"b70700f0",
         369 => x"03a54702",
         370 => x"13754500",
         371 => x"67800000",
         372 => x"370700f0",
         373 => x"13070702",
         374 => x"83274700",
         375 => x"93f74700",
         376 => x"e38c07fe",
         377 => x"03258700",
         378 => x"1375f50f",
         379 => x"67800000",
         380 => x"130101fd",
         381 => x"232e3101",
         382 => x"b7190010",
         383 => x"23248102",
         384 => x"23229102",
         385 => x"23202103",
         386 => x"232c4101",
         387 => x"232a5101",
         388 => x"23286101",
         389 => x"23267101",
         390 => x"23261102",
         391 => x"93040500",
         392 => x"13040000",
         393 => x"9389c9b5",
         394 => x"13095001",
         395 => x"138bf5ff",
         396 => x"130a2000",
         397 => x"930a2001",
         398 => x"b71b0010",
         399 => x"eff05ff9",
         400 => x"1377f50f",
         401 => x"6340e902",
         402 => x"6352ea02",
         403 => x"9307d7ff",
         404 => x"63eefa00",
         405 => x"93972700",
         406 => x"b387f900",
         407 => x"83a70700",
         408 => x"67800700",
         409 => x"9307f007",
         410 => x"630cf706",
         411 => x"6352640f",
         412 => x"9377f50f",
         413 => x"938607fe",
         414 => x"93f6f60f",
         415 => x"1306e005",
         416 => x"e36ed6fa",
         417 => x"b3868400",
         418 => x"2380f600",
         419 => x"13050700",
         420 => x"13041400",
         421 => x"ef008011",
         422 => x"6ff05ffa",
         423 => x"b3848400",
         424 => x"37150010",
         425 => x"23800400",
         426 => x"130585cd",
         427 => x"ef000012",
         428 => x"8320c102",
         429 => x"13050400",
         430 => x"03248102",
         431 => x"83244102",
         432 => x"03290102",
         433 => x"8329c101",
         434 => x"032a8101",
         435 => x"832a4101",
         436 => x"032b0101",
         437 => x"832bc100",
         438 => x"13010103",
         439 => x"67800000",
         440 => x"635a8002",
         441 => x"1305f007",
         442 => x"ef00400c",
         443 => x"1304f4ff",
         444 => x"6ff0dff4",
         445 => x"1385cbca",
         446 => x"ef00400d",
         447 => x"eff05fed",
         448 => x"1377f50f",
         449 => x"13040000",
         450 => x"e350e9f4",
         451 => x"9307f007",
         452 => x"e31ef7f4",
         453 => x"23248101",
         454 => x"130c5001",
         455 => x"13057000",
         456 => x"ef00c008",
         457 => x"eff0dfea",
         458 => x"1377f50f",
         459 => x"6348ec02",
         460 => x"032c8100",
         461 => x"6ff05ff1",
         462 => x"635a8002",
         463 => x"1305f007",
         464 => x"1304f4ff",
         465 => x"ef008006",
         466 => x"e31a04fe",
         467 => x"6ff01fef",
         468 => x"13057000",
         469 => x"ef008005",
         470 => x"6ff05fee",
         471 => x"9307f007",
         472 => x"e30ef7fa",
         473 => x"032c8100",
         474 => x"6ff05ff0",
         475 => x"eff05fe6",
         476 => x"1377f50f",
         477 => x"93075001",
         478 => x"e3d8e7ec",
         479 => x"6ff01ff9",
         480 => x"f32710fc",
         481 => x"63960700",
         482 => x"b7f7fa02",
         483 => x"93870708",
         484 => x"63060500",
         485 => x"33d5a702",
         486 => x"1305f5ff",
         487 => x"b70700f0",
         488 => x"23a6a702",
         489 => x"23a0b702",
         490 => x"67800000",
         491 => x"370700f0",
         492 => x"1375f50f",
         493 => x"13070702",
         494 => x"2324a700",
         495 => x"83274700",
         496 => x"93f70701",
         497 => x"e38c07fe",
         498 => x"67800000",
         499 => x"630e0502",
         500 => x"130101ff",
         501 => x"23248100",
         502 => x"23261100",
         503 => x"13040500",
         504 => x"03450500",
         505 => x"630a0500",
         506 => x"13041400",
         507 => x"eff01ffc",
         508 => x"03450400",
         509 => x"e31a05fe",
         510 => x"8320c100",
         511 => x"03248100",
         512 => x"13010101",
         513 => x"67800000",
         514 => x"67800000",
         515 => x"130101fe",
         516 => x"232e1100",
         517 => x"232c8100",
         518 => x"6350a00a",
         519 => x"23263101",
         520 => x"b7190010",
         521 => x"232a9100",
         522 => x"23282101",
         523 => x"23244101",
         524 => x"13090500",
         525 => x"93040000",
         526 => x"13040000",
         527 => x"938999ba",
         528 => x"130a1000",
         529 => x"6f000001",
         530 => x"3364c400",
         531 => x"93841400",
         532 => x"63029904",
         533 => x"eff0dfd7",
         534 => x"b387a900",
         535 => x"83c70700",
         536 => x"130605fd",
         537 => x"13144400",
         538 => x"13f74700",
         539 => x"93f64704",
         540 => x"e31c07fc",
         541 => x"93f73700",
         542 => x"e38a06fc",
         543 => x"63944701",
         544 => x"13050502",
         545 => x"130595fa",
         546 => x"93841400",
         547 => x"3364a400",
         548 => x"e31299fc",
         549 => x"8320c101",
         550 => x"13050400",
         551 => x"03248101",
         552 => x"83244101",
         553 => x"03290101",
         554 => x"8329c100",
         555 => x"032a8100",
         556 => x"13010102",
         557 => x"67800000",
         558 => x"13040000",
         559 => x"8320c101",
         560 => x"13050400",
         561 => x"03248101",
         562 => x"13010102",
         563 => x"67800000",
         564 => x"83470500",
         565 => x"37160010",
         566 => x"130696ba",
         567 => x"3307f600",
         568 => x"03470700",
         569 => x"93060500",
         570 => x"13758700",
         571 => x"630e0500",
         572 => x"83c71600",
         573 => x"93861600",
         574 => x"3307f600",
         575 => x"03470700",
         576 => x"13758700",
         577 => x"e31605fe",
         578 => x"13754704",
         579 => x"630a0506",
         580 => x"13050000",
         581 => x"13031000",
         582 => x"6f000002",
         583 => x"83c71600",
         584 => x"33e5a800",
         585 => x"93861600",
         586 => x"3307f600",
         587 => x"03470700",
         588 => x"13784704",
         589 => x"63000804",
         590 => x"13784700",
         591 => x"938807fd",
         592 => x"13773700",
         593 => x"13154500",
         594 => x"e31a08fc",
         595 => x"63146700",
         596 => x"93870702",
         597 => x"938797fa",
         598 => x"33e5a700",
         599 => x"83c71600",
         600 => x"93861600",
         601 => x"3307f600",
         602 => x"03470700",
         603 => x"13784704",
         604 => x"e31408fc",
         605 => x"63840500",
         606 => x"23a0d500",
         607 => x"67800000",
         608 => x"13050000",
         609 => x"6ff01fff",
         610 => x"130101fe",
         611 => x"232e1100",
         612 => x"23220100",
         613 => x"23240100",
         614 => x"23260100",
         615 => x"63040506",
         616 => x"232c8100",
         617 => x"93070500",
         618 => x"13040500",
         619 => x"63440504",
         620 => x"13074100",
         621 => x"1306a000",
         622 => x"13089000",
         623 => x"b3f6c702",
         624 => x"13050700",
         625 => x"1307f7ff",
         626 => x"93850700",
         627 => x"93860603",
         628 => x"a305d700",
         629 => x"b3d7c702",
         630 => x"e362b8fe",
         631 => x"3305c500",
         632 => x"eff0dfde",
         633 => x"8320c101",
         634 => x"03248101",
         635 => x"13010102",
         636 => x"67800000",
         637 => x"1305d002",
         638 => x"eff05fdb",
         639 => x"b3078040",
         640 => x"6ff01ffb",
         641 => x"13050003",
         642 => x"eff05fda",
         643 => x"8320c101",
         644 => x"13010102",
         645 => x"67800000",
         646 => x"130101fe",
         647 => x"232e1100",
         648 => x"23220100",
         649 => x"23240100",
         650 => x"23060100",
         651 => x"9387f5ff",
         652 => x"13077000",
         653 => x"6376f700",
         654 => x"93077000",
         655 => x"93058000",
         656 => x"13074100",
         657 => x"b307f700",
         658 => x"b385b740",
         659 => x"13069003",
         660 => x"9376f500",
         661 => x"13870603",
         662 => x"6374e600",
         663 => x"13877605",
         664 => x"2380e700",
         665 => x"9387f7ff",
         666 => x"13554500",
         667 => x"e392f5fe",
         668 => x"13054100",
         669 => x"eff09fd5",
         670 => x"8320c101",
         671 => x"13010102",
         672 => x"67800000",
         673 => x"130101ff",
         674 => x"23248100",
         675 => x"23229100",
         676 => x"37140010",
         677 => x"b7140010",
         678 => x"9387c4e1",
         679 => x"1304c4e1",
         680 => x"3304f440",
         681 => x"23202101",
         682 => x"23261100",
         683 => x"13542440",
         684 => x"9384c4e1",
         685 => x"13090000",
         686 => x"63108904",
         687 => x"b7140010",
         688 => x"37140010",
         689 => x"9387c4e1",
         690 => x"1304c4e1",
         691 => x"3304f440",
         692 => x"13542440",
         693 => x"9384c4e1",
         694 => x"13090000",
         695 => x"63188902",
         696 => x"8320c100",
         697 => x"03248100",
         698 => x"83244100",
         699 => x"03290100",
         700 => x"13010101",
         701 => x"67800000",
         702 => x"83a70400",
         703 => x"13091900",
         704 => x"93844400",
         705 => x"e7800700",
         706 => x"6ff01ffb",
         707 => x"83a70400",
         708 => x"13091900",
         709 => x"93844400",
         710 => x"e7800700",
         711 => x"6ff01ffc",
         712 => x"630a0602",
         713 => x"1306f6ff",
         714 => x"13070000",
         715 => x"b307e500",
         716 => x"b386e500",
         717 => x"83c70700",
         718 => x"83c60600",
         719 => x"6398d700",
         720 => x"6306c700",
         721 => x"13071700",
         722 => x"e39207fe",
         723 => x"3385d740",
         724 => x"67800000",
         725 => x"13050000",
         726 => x"67800000",
         727 => x"f4060010",
         728 => x"6c060010",
         729 => x"6c060010",
         730 => x"6c060010",
         731 => x"6c060010",
         732 => x"e0060010",
         733 => x"6c060010",
         734 => x"9c060010",
         735 => x"6c060010",
         736 => x"6c060010",
         737 => x"9c060010",
         738 => x"6c060010",
         739 => x"6c060010",
         740 => x"6c060010",
         741 => x"6c060010",
         742 => x"6c060010",
         743 => x"6c060010",
         744 => x"6c060010",
         745 => x"38070010",
         746 => x"00202020",
         747 => x"20202020",
         748 => x"20202828",
         749 => x"28282820",
         750 => x"20202020",
         751 => x"20202020",
         752 => x"20202020",
         753 => x"20202020",
         754 => x"20881010",
         755 => x"10101010",
         756 => x"10101010",
         757 => x"10101010",
         758 => x"10040404",
         759 => x"04040404",
         760 => x"04040410",
         761 => x"10101010",
         762 => x"10104141",
         763 => x"41414141",
         764 => x"01010101",
         765 => x"01010101",
         766 => x"01010101",
         767 => x"01010101",
         768 => x"01010101",
         769 => x"10101010",
         770 => x"10104242",
         771 => x"42424242",
         772 => x"02020202",
         773 => x"02020202",
         774 => x"02020202",
         775 => x"02020202",
         776 => x"02020202",
         777 => x"10101010",
         778 => x"20000000",
         779 => x"00000000",
         780 => x"00000000",
         781 => x"00000000",
         782 => x"00000000",
         783 => x"00000000",
         784 => x"00000000",
         785 => x"00000000",
         786 => x"00000000",
         787 => x"00000000",
         788 => x"00000000",
         789 => x"00000000",
         790 => x"00000000",
         791 => x"00000000",
         792 => x"00000000",
         793 => x"00000000",
         794 => x"00000000",
         795 => x"00000000",
         796 => x"00000000",
         797 => x"00000000",
         798 => x"00000000",
         799 => x"00000000",
         800 => x"00000000",
         801 => x"00000000",
         802 => x"00000000",
         803 => x"00000000",
         804 => x"00000000",
         805 => x"00000000",
         806 => x"00000000",
         807 => x"00000000",
         808 => x"00000000",
         809 => x"00000000",
         810 => x"00000000",
         811 => x"3c627265",
         812 => x"616b3e0d",
         813 => x"0a000000",
         814 => x"0d0a5448",
         815 => x"55415320",
         816 => x"52495343",
         817 => x"2d562042",
         818 => x"6f6f746c",
         819 => x"6f616465",
         820 => x"72207630",
         821 => x"2e352e31",
         822 => x"0d0a0000",
         823 => x"436c6f63",
         824 => x"6b206672",
         825 => x"65717565",
         826 => x"6e63793a",
         827 => x"20000000",
         828 => x"3f0a0000",
         829 => x"3e200000",
         830 => x"68000000",
         831 => x"48656c70",
         832 => x"3a0d0a20",
         833 => x"68202020",
         834 => x"20202020",
         835 => x"20202020",
         836 => x"20202020",
         837 => x"202d2074",
         838 => x"68697320",
         839 => x"68656c70",
         840 => x"0d0a2072",
         841 => x"20202020",
         842 => x"20202020",
         843 => x"20202020",
         844 => x"20202020",
         845 => x"2d207275",
         846 => x"6e206170",
         847 => x"706c6963",
         848 => x"6174696f",
         849 => x"6e0d0a20",
         850 => x"7277203c",
         851 => x"61646472",
         852 => x"3e202020",
         853 => x"20202020",
         854 => x"202d2072",
         855 => x"65616420",
         856 => x"776f7264",
         857 => x"2066726f",
         858 => x"6d206164",
         859 => x"64720d0a",
         860 => x"20777720",
         861 => x"3c616464",
         862 => x"723e203c",
         863 => x"64617461",
         864 => x"3e202d20",
         865 => x"77726974",
         866 => x"6520776f",
         867 => x"72642064",
         868 => x"61746120",
         869 => x"61742061",
         870 => x"6464720d",
         871 => x"0a206477",
         872 => x"203c6164",
         873 => x"64723e20",
         874 => x"20202020",
         875 => x"2020202d",
         876 => x"2064756d",
         877 => x"70203136",
         878 => x"20776f72",
         879 => x"64730d0a",
         880 => x"206e2020",
         881 => x"20202020",
         882 => x"20202020",
         883 => x"20202020",
         884 => x"20202d20",
         885 => x"64756d70",
         886 => x"206e6578",
         887 => x"74203136",
         888 => x"20776f72",
         889 => x"64730000",
         890 => x"72000000",
         891 => x"72772000",
         892 => x"3a200000",
         893 => x"4e6f7420",
         894 => x"6f6e2034",
         895 => x"2d627974",
         896 => x"6520626f",
         897 => x"756e6461",
         898 => x"72792100",
         899 => x"77772000",
         900 => x"64772000",
         901 => x"20200000",
         902 => x"3f3f0000",
         903 => x"00000000"
            );
end package bootrom_image;
