-- srec2vhdl table generator
-- for input file 'bootloader.srec'
-- date: Sun Nov 19 13:42:45 2023


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package bootrom_image is
    constant bootrom_contents : memory_type := (
           0 => x"97020000",
           1 => x"93824256",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"b7070020",
           9 => x"93870700",
          10 => x"13070500",
          11 => x"3386e740",
          12 => x"63f4e700",
          13 => x"13060000",
          14 => x"93050000",
          15 => x"13050500",
          16 => x"ef008052",
          17 => x"37050020",
          18 => x"b7070020",
          19 => x"93870700",
          20 => x"13070500",
          21 => x"3386e740",
          22 => x"63f4e700",
          23 => x"13060000",
          24 => x"b7150010",
          25 => x"938545e4",
          26 => x"13050500",
          27 => x"ef008051",
          28 => x"ef00d021",
          29 => x"37c50100",
          30 => x"93050000",
          31 => x"13050520",
          32 => x"ef008070",
          33 => x"37150010",
          34 => x"130505ce",
          35 => x"ef008074",
          36 => x"37150010",
          37 => x"130545d0",
          38 => x"ef00c073",
          39 => x"732510fc",
          40 => x"37190010",
          41 => x"ef00d00e",
          42 => x"130509cd",
          43 => x"ef008072",
          44 => x"b70700f0",
          45 => x"1307f03f",
          46 => x"370a1000",
          47 => x"b709a000",
          48 => x"23a2e700",
          49 => x"93041000",
          50 => x"130afaff",
          51 => x"b70a00f0",
          52 => x"93891900",
          53 => x"b3f74401",
          54 => x"639c0700",
          55 => x"1305a002",
          56 => x"ef00406d",
          57 => x"83a74a00",
          58 => x"93d71700",
          59 => x"23a2fa00",
          60 => x"ef00804d",
          61 => x"13040500",
          62 => x"63160504",
          63 => x"93841400",
          64 => x"e39a34fd",
          65 => x"b70700f0",
          66 => x"23a20700",
          67 => x"631a0400",
          68 => x"93050000",
          69 => x"13050000",
          70 => x"ef000067",
          71 => x"e7000400",
          72 => x"ef00804b",
          73 => x"1375f50f",
          74 => x"93071002",
          75 => x"6300f502",
          76 => x"93074002",
          77 => x"93040000",
          78 => x"6316f520",
          79 => x"13041000",
          80 => x"6f00c001",
          81 => x"13041000",
          82 => x"6ff0dffb",
          83 => x"37150010",
          84 => x"130585d1",
          85 => x"ef000068",
          86 => x"13040000",
          87 => x"93040000",
          88 => x"370a00f0",
          89 => x"130b3005",
          90 => x"930ba004",
          91 => x"130c3002",
          92 => x"93092000",
          93 => x"930ca000",
          94 => x"b71a0010",
          95 => x"83274a00",
          96 => x"93c71700",
          97 => x"2322fa00",
          98 => x"ef000045",
          99 => x"1375f50f",
         100 => x"631e6517",
         101 => x"ef004044",
         102 => x"137df50f",
         103 => x"9307fdfc",
         104 => x"93f7f70f",
         105 => x"63e6f910",
         106 => x"93071003",
         107 => x"631afd04",
         108 => x"13052000",
         109 => x"ef000066",
         110 => x"930dd5ff",
         111 => x"13054000",
         112 => x"ef004065",
         113 => x"b70601ff",
         114 => x"b705ffff",
         115 => x"130d0500",
         116 => x"b38dad00",
         117 => x"9386f6ff",
         118 => x"9385f50f",
         119 => x"6398ad05",
         120 => x"130da000",
         121 => x"ef00403f",
         122 => x"1375f50f",
         123 => x"e31ca5ff",
         124 => x"e31604f8",
         125 => x"13858ad1",
         126 => x"ef00c05d",
         127 => x"6ff01ff8",
         128 => x"93072003",
         129 => x"13052000",
         130 => x"631afd00",
         131 => x"ef008060",
         132 => x"930dc5ff",
         133 => x"13056000",
         134 => x"6ff09ffa",
         135 => x"ef00805f",
         136 => x"930db5ff",
         137 => x"13058000",
         138 => x"6ff09ff9",
         139 => x"1378cdff",
         140 => x"13052000",
         141 => x"2326b100",
         142 => x"2324d100",
         143 => x"23220101",
         144 => x"ef00405d",
         145 => x"03284100",
         146 => x"93070500",
         147 => x"37060001",
         148 => x"13753d00",
         149 => x"03270800",
         150 => x"83268100",
         151 => x"8325c100",
         152 => x"93083000",
         153 => x"1306f6ff",
         154 => x"13031000",
         155 => x"63063503",
         156 => x"630a1503",
         157 => x"630c6500",
         158 => x"137707f0",
         159 => x"b3e7e700",
         160 => x"2320f800",
         161 => x"130d1d00",
         162 => x"6ff05ff5",
         163 => x"3377b700",
         164 => x"93978700",
         165 => x"6ff09ffe",
         166 => x"3377d700",
         167 => x"93970701",
         168 => x"6ff0dffd",
         169 => x"3377c700",
         170 => x"93978701",
         171 => x"6ff01ffd",
         172 => x"93079dfc",
         173 => x"93f7f70f",
         174 => x"63e2f904",
         175 => x"13052000",
         176 => x"ef004055",
         177 => x"93077003",
         178 => x"13058000",
         179 => x"630afd00",
         180 => x"93078003",
         181 => x"13056000",
         182 => x"6304fd00",
         183 => x"13054000",
         184 => x"ef004053",
         185 => x"93040500",
         186 => x"130da000",
         187 => x"ef00c02e",
         188 => x"1375f50f",
         189 => x"e31ca5ff",
         190 => x"6ff09fef",
         191 => x"ef00c02d",
         192 => x"1375f50f",
         193 => x"e31c95ff",
         194 => x"6ff09fee",
         195 => x"631c7509",
         196 => x"63180400",
         197 => x"37150010",
         198 => x"130585d1",
         199 => x"ef00804b",
         200 => x"93050000",
         201 => x"13050000",
         202 => x"ef000046",
         203 => x"b70700f0",
         204 => x"23a20700",
         205 => x"e7800400",
         206 => x"b70700f0",
         207 => x"1307a00a",
         208 => x"23a2e700",
         209 => x"130509cd",
         210 => x"b7190010",
         211 => x"ef008048",
         212 => x"13040000",
         213 => x"b71b0010",
         214 => x"9389d9bc",
         215 => x"b7170010",
         216 => x"1385c7d1",
         217 => x"ef000047",
         218 => x"93059002",
         219 => x"13054101",
         220 => x"ef008028",
         221 => x"13054101",
         222 => x"ef00c07e",
         223 => x"b7170010",
         224 => x"130a0500",
         225 => x"938507d2",
         226 => x"13054101",
         227 => x"ef00c021",
         228 => x"631e0500",
         229 => x"37150010",
         230 => x"130545d2",
         231 => x"ef008043",
         232 => x"6f004003",
         233 => x"e31685e5",
         234 => x"6ff01ff9",
         235 => x"b7170010",
         236 => x"938507e1",
         237 => x"13054101",
         238 => x"ef00001f",
         239 => x"63100502",
         240 => x"93050000",
         241 => x"ef00403c",
         242 => x"b70700f0",
         243 => x"23a20700",
         244 => x"e7800400",
         245 => x"e3040af8",
         246 => x"6f000018",
         247 => x"b7170010",
         248 => x"13063000",
         249 => x"938547e1",
         250 => x"13054101",
         251 => x"ef00c073",
         252 => x"63100504",
         253 => x"93050000",
         254 => x"13057101",
         255 => x"ef00c04d",
         256 => x"93773500",
         257 => x"13040500",
         258 => x"63960706",
         259 => x"93058000",
         260 => x"ef000061",
         261 => x"37150010",
         262 => x"130585e1",
         263 => x"ef00803b",
         264 => x"03250400",
         265 => x"93058000",
         266 => x"ef00805f",
         267 => x"6ff09ffa",
         268 => x"b7170010",
         269 => x"13063000",
         270 => x"938547e3",
         271 => x"13054101",
         272 => x"ef00806e",
         273 => x"631e0502",
         274 => x"93050101",
         275 => x"13057101",
         276 => x"ef008048",
         277 => x"93773500",
         278 => x"13040500",
         279 => x"639c0700",
         280 => x"03250101",
         281 => x"93050000",
         282 => x"ef000047",
         283 => x"2320a400",
         284 => x"6ff05ff6",
         285 => x"37150010",
         286 => x"1305c5e1",
         287 => x"6ff01ff2",
         288 => x"13063000",
         289 => x"93858be3",
         290 => x"13054101",
         291 => x"ef00c069",
         292 => x"83474101",
         293 => x"1307e006",
         294 => x"63080508",
         295 => x"6396e70a",
         296 => x"93773400",
         297 => x"e39807fc",
         298 => x"130c0404",
         299 => x"b71c0010",
         300 => x"371d0010",
         301 => x"930d80ff",
         302 => x"93058000",
         303 => x"13050400",
         304 => x"ef000056",
         305 => x"13858ce1",
         306 => x"ef00c030",
         307 => x"032a0400",
         308 => x"93058000",
         309 => x"930a8001",
         310 => x"13050a00",
         311 => x"ef004054",
         312 => x"1305cde3",
         313 => x"ef00002f",
         314 => x"370b00ff",
         315 => x"33756a01",
         316 => x"33555501",
         317 => x"b3063501",
         318 => x"83c60600",
         319 => x"93f67609",
         320 => x"63800604",
         321 => x"938a8aff",
         322 => x"ef00c02a",
         323 => x"135b8b00",
         324 => x"e39ebafd",
         325 => x"13044400",
         326 => x"130509cd",
         327 => x"ef00802b",
         328 => x"e31c8cf8",
         329 => x"6ff09fe3",
         330 => x"e38ce7f6",
         331 => x"93050000",
         332 => x"13057101",
         333 => x"ef00403a",
         334 => x"13040500",
         335 => x"6ff05ff6",
         336 => x"1305e002",
         337 => x"6ff01ffc",
         338 => x"e30a0ae0",
         339 => x"37150010",
         340 => x"130505e4",
         341 => x"ef000028",
         342 => x"130509cd",
         343 => x"ef008027",
         344 => x"6ff0dfdf",
         345 => x"6f000000",
         346 => x"13030500",
         347 => x"630a0600",
         348 => x"2300b300",
         349 => x"1306f6ff",
         350 => x"13031300",
         351 => x"e31a06fe",
         352 => x"67800000",
         353 => x"13030500",
         354 => x"630e0600",
         355 => x"83830500",
         356 => x"23007300",
         357 => x"1306f6ff",
         358 => x"13031300",
         359 => x"93851500",
         360 => x"e31606fe",
         361 => x"67800000",
         362 => x"03460500",
         363 => x"83c60500",
         364 => x"13051500",
         365 => x"93851500",
         366 => x"6314d600",
         367 => x"e31606fe",
         368 => x"3305d640",
         369 => x"67800000",
         370 => x"b70700f0",
         371 => x"03a54702",
         372 => x"13754500",
         373 => x"67800000",
         374 => x"370700f0",
         375 => x"13070702",
         376 => x"83274700",
         377 => x"93f74700",
         378 => x"e38c07fe",
         379 => x"03258700",
         380 => x"1375f50f",
         381 => x"67800000",
         382 => x"130101fd",
         383 => x"232e3101",
         384 => x"b7190010",
         385 => x"23248102",
         386 => x"23229102",
         387 => x"23202103",
         388 => x"232c4101",
         389 => x"232a5101",
         390 => x"23286101",
         391 => x"23267101",
         392 => x"23261102",
         393 => x"93040500",
         394 => x"13040000",
         395 => x"938909b8",
         396 => x"13095001",
         397 => x"138bf5ff",
         398 => x"130a2000",
         399 => x"930a2001",
         400 => x"b71b0010",
         401 => x"eff05ff9",
         402 => x"1377f50f",
         403 => x"6340e902",
         404 => x"6352ea02",
         405 => x"9307d7ff",
         406 => x"63eefa00",
         407 => x"93972700",
         408 => x"b387f900",
         409 => x"83a70700",
         410 => x"67800700",
         411 => x"9307f007",
         412 => x"630cf706",
         413 => x"6352640f",
         414 => x"9377f50f",
         415 => x"938607fe",
         416 => x"93f6f60f",
         417 => x"1306e005",
         418 => x"e36ed6fa",
         419 => x"b3868400",
         420 => x"2380f600",
         421 => x"13050700",
         422 => x"13041400",
         423 => x"ef008011",
         424 => x"6ff05ffa",
         425 => x"b3848400",
         426 => x"37150010",
         427 => x"23800400",
         428 => x"130505cd",
         429 => x"ef000012",
         430 => x"8320c102",
         431 => x"13050400",
         432 => x"03248102",
         433 => x"83244102",
         434 => x"03290102",
         435 => x"8329c101",
         436 => x"032a8101",
         437 => x"832a4101",
         438 => x"032b0101",
         439 => x"832bc100",
         440 => x"13010103",
         441 => x"67800000",
         442 => x"635a8002",
         443 => x"1305f007",
         444 => x"ef00400c",
         445 => x"1304f4ff",
         446 => x"6ff0dff4",
         447 => x"13854bcd",
         448 => x"ef00400d",
         449 => x"eff05fed",
         450 => x"1377f50f",
         451 => x"13040000",
         452 => x"e350e9f4",
         453 => x"9307f007",
         454 => x"e31ef7f4",
         455 => x"23248101",
         456 => x"130c5001",
         457 => x"13057000",
         458 => x"ef00c008",
         459 => x"eff0dfea",
         460 => x"1377f50f",
         461 => x"6348ec02",
         462 => x"032c8100",
         463 => x"6ff05ff1",
         464 => x"635a8002",
         465 => x"1305f007",
         466 => x"1304f4ff",
         467 => x"ef008006",
         468 => x"e31a04fe",
         469 => x"6ff01fef",
         470 => x"13057000",
         471 => x"ef008005",
         472 => x"6ff05fee",
         473 => x"9307f007",
         474 => x"e30ef7fa",
         475 => x"032c8100",
         476 => x"6ff05ff0",
         477 => x"eff05fe6",
         478 => x"1377f50f",
         479 => x"93075001",
         480 => x"e3d8e7ec",
         481 => x"6ff01ff9",
         482 => x"f32710fc",
         483 => x"63960700",
         484 => x"b7f7fa02",
         485 => x"93870708",
         486 => x"63060500",
         487 => x"33d5a702",
         488 => x"1305f5ff",
         489 => x"b70700f0",
         490 => x"23a6a702",
         491 => x"23a0b702",
         492 => x"67800000",
         493 => x"370700f0",
         494 => x"1375f50f",
         495 => x"13070702",
         496 => x"2324a700",
         497 => x"83274700",
         498 => x"93f70701",
         499 => x"e38c07fe",
         500 => x"67800000",
         501 => x"630e0502",
         502 => x"130101ff",
         503 => x"23248100",
         504 => x"23261100",
         505 => x"13040500",
         506 => x"03450500",
         507 => x"630a0500",
         508 => x"13041400",
         509 => x"eff01ffc",
         510 => x"03450400",
         511 => x"e31a05fe",
         512 => x"8320c100",
         513 => x"03248100",
         514 => x"13010101",
         515 => x"67800000",
         516 => x"67800000",
         517 => x"130101fe",
         518 => x"232e1100",
         519 => x"232c8100",
         520 => x"6350a00a",
         521 => x"23263101",
         522 => x"b7190010",
         523 => x"232a9100",
         524 => x"23282101",
         525 => x"23244101",
         526 => x"13090500",
         527 => x"93040000",
         528 => x"13040000",
         529 => x"9389d9bc",
         530 => x"130a1000",
         531 => x"6f000001",
         532 => x"3364c400",
         533 => x"93841400",
         534 => x"63029904",
         535 => x"eff0dfd7",
         536 => x"b387a900",
         537 => x"83c70700",
         538 => x"130605fd",
         539 => x"13144400",
         540 => x"13f74700",
         541 => x"93f64704",
         542 => x"e31c07fc",
         543 => x"93f73700",
         544 => x"e38a06fc",
         545 => x"63944701",
         546 => x"13050502",
         547 => x"130595fa",
         548 => x"93841400",
         549 => x"3364a400",
         550 => x"e31299fc",
         551 => x"8320c101",
         552 => x"13050400",
         553 => x"03248101",
         554 => x"83244101",
         555 => x"03290101",
         556 => x"8329c100",
         557 => x"032a8100",
         558 => x"13010102",
         559 => x"67800000",
         560 => x"13040000",
         561 => x"8320c101",
         562 => x"13050400",
         563 => x"03248101",
         564 => x"13010102",
         565 => x"67800000",
         566 => x"83470500",
         567 => x"37160010",
         568 => x"1306d6bc",
         569 => x"3307f600",
         570 => x"03470700",
         571 => x"93060500",
         572 => x"13758700",
         573 => x"630e0500",
         574 => x"83c71600",
         575 => x"93861600",
         576 => x"3307f600",
         577 => x"03470700",
         578 => x"13758700",
         579 => x"e31605fe",
         580 => x"13754704",
         581 => x"630a0506",
         582 => x"13050000",
         583 => x"13031000",
         584 => x"6f000002",
         585 => x"83c71600",
         586 => x"33e5a800",
         587 => x"93861600",
         588 => x"3307f600",
         589 => x"03470700",
         590 => x"13784704",
         591 => x"63000804",
         592 => x"13784700",
         593 => x"938807fd",
         594 => x"13773700",
         595 => x"13154500",
         596 => x"e31a08fc",
         597 => x"63146700",
         598 => x"93870702",
         599 => x"938797fa",
         600 => x"33e5a700",
         601 => x"83c71600",
         602 => x"93861600",
         603 => x"3307f600",
         604 => x"03470700",
         605 => x"13784704",
         606 => x"e31408fc",
         607 => x"63840500",
         608 => x"23a0d500",
         609 => x"67800000",
         610 => x"13050000",
         611 => x"6ff01fff",
         612 => x"130101fe",
         613 => x"232e1100",
         614 => x"23220100",
         615 => x"23240100",
         616 => x"23260100",
         617 => x"63040506",
         618 => x"232c8100",
         619 => x"93070500",
         620 => x"13040500",
         621 => x"63440504",
         622 => x"13074100",
         623 => x"1306a000",
         624 => x"13089000",
         625 => x"b3f6c702",
         626 => x"13050700",
         627 => x"1307f7ff",
         628 => x"93850700",
         629 => x"93860603",
         630 => x"a305d700",
         631 => x"b3d7c702",
         632 => x"e362b8fe",
         633 => x"3305c500",
         634 => x"eff0dfde",
         635 => x"8320c101",
         636 => x"03248101",
         637 => x"13010102",
         638 => x"67800000",
         639 => x"1305d002",
         640 => x"eff05fdb",
         641 => x"b3078040",
         642 => x"6ff01ffb",
         643 => x"13050003",
         644 => x"eff05fda",
         645 => x"8320c101",
         646 => x"13010102",
         647 => x"67800000",
         648 => x"130101fe",
         649 => x"232e1100",
         650 => x"23220100",
         651 => x"23240100",
         652 => x"23060100",
         653 => x"9387f5ff",
         654 => x"13077000",
         655 => x"6376f700",
         656 => x"93077000",
         657 => x"93058000",
         658 => x"13074100",
         659 => x"b307f700",
         660 => x"b385b740",
         661 => x"13069003",
         662 => x"9376f500",
         663 => x"13870603",
         664 => x"6374e600",
         665 => x"13877605",
         666 => x"2380e700",
         667 => x"9387f7ff",
         668 => x"13554500",
         669 => x"e392f5fe",
         670 => x"13054100",
         671 => x"eff09fd5",
         672 => x"8320c101",
         673 => x"13010102",
         674 => x"67800000",
         675 => x"130101ff",
         676 => x"23248100",
         677 => x"23229100",
         678 => x"37140010",
         679 => x"b7140010",
         680 => x"938744e4",
         681 => x"130444e4",
         682 => x"3304f440",
         683 => x"23202101",
         684 => x"23261100",
         685 => x"13542440",
         686 => x"938444e4",
         687 => x"13090000",
         688 => x"63108904",
         689 => x"b7140010",
         690 => x"37140010",
         691 => x"938744e4",
         692 => x"130444e4",
         693 => x"3304f440",
         694 => x"13542440",
         695 => x"938444e4",
         696 => x"13090000",
         697 => x"63188902",
         698 => x"8320c100",
         699 => x"03248100",
         700 => x"83244100",
         701 => x"03290100",
         702 => x"13010101",
         703 => x"67800000",
         704 => x"83a70400",
         705 => x"13091900",
         706 => x"93844400",
         707 => x"e7800700",
         708 => x"6ff01ffb",
         709 => x"83a70400",
         710 => x"13091900",
         711 => x"93844400",
         712 => x"e7800700",
         713 => x"6ff01ffc",
         714 => x"630a0602",
         715 => x"1306f6ff",
         716 => x"13070000",
         717 => x"b307e500",
         718 => x"b386e500",
         719 => x"83c70700",
         720 => x"83c60600",
         721 => x"6398d700",
         722 => x"6306c700",
         723 => x"13071700",
         724 => x"e39207fe",
         725 => x"3385d740",
         726 => x"67800000",
         727 => x"13050000",
         728 => x"67800000",
         729 => x"93070500",
         730 => x"03c70700",
         731 => x"93871700",
         732 => x"e31c07fe",
         733 => x"3385a740",
         734 => x"1305f5ff",
         735 => x"67800000",
         736 => x"fc060010",
         737 => x"74060010",
         738 => x"74060010",
         739 => x"74060010",
         740 => x"74060010",
         741 => x"e8060010",
         742 => x"74060010",
         743 => x"a4060010",
         744 => x"74060010",
         745 => x"74060010",
         746 => x"a4060010",
         747 => x"74060010",
         748 => x"74060010",
         749 => x"74060010",
         750 => x"74060010",
         751 => x"74060010",
         752 => x"74060010",
         753 => x"74060010",
         754 => x"40070010",
         755 => x"00202020",
         756 => x"20202020",
         757 => x"20202828",
         758 => x"28282820",
         759 => x"20202020",
         760 => x"20202020",
         761 => x"20202020",
         762 => x"20202020",
         763 => x"20881010",
         764 => x"10101010",
         765 => x"10101010",
         766 => x"10101010",
         767 => x"10040404",
         768 => x"04040404",
         769 => x"04040410",
         770 => x"10101010",
         771 => x"10104141",
         772 => x"41414141",
         773 => x"01010101",
         774 => x"01010101",
         775 => x"01010101",
         776 => x"01010101",
         777 => x"01010101",
         778 => x"10101010",
         779 => x"10104242",
         780 => x"42424242",
         781 => x"02020202",
         782 => x"02020202",
         783 => x"02020202",
         784 => x"02020202",
         785 => x"02020202",
         786 => x"10101010",
         787 => x"20000000",
         788 => x"00000000",
         789 => x"00000000",
         790 => x"00000000",
         791 => x"00000000",
         792 => x"00000000",
         793 => x"00000000",
         794 => x"00000000",
         795 => x"00000000",
         796 => x"00000000",
         797 => x"00000000",
         798 => x"00000000",
         799 => x"00000000",
         800 => x"00000000",
         801 => x"00000000",
         802 => x"00000000",
         803 => x"00000000",
         804 => x"00000000",
         805 => x"00000000",
         806 => x"00000000",
         807 => x"00000000",
         808 => x"00000000",
         809 => x"00000000",
         810 => x"00000000",
         811 => x"00000000",
         812 => x"00000000",
         813 => x"00000000",
         814 => x"00000000",
         815 => x"00000000",
         816 => x"00000000",
         817 => x"00000000",
         818 => x"00000000",
         819 => x"00000000",
         820 => x"0d0a0000",
         821 => x"3c627265",
         822 => x"616b3e0d",
         823 => x"0a000000",
         824 => x"0d0a5448",
         825 => x"55415320",
         826 => x"52495343",
         827 => x"2d562042",
         828 => x"6f6f746c",
         829 => x"6f616465",
         830 => x"72207630",
         831 => x"2e350d0a",
         832 => x"00000000",
         833 => x"436c6f63",
         834 => x"6b206672",
         835 => x"65717565",
         836 => x"6e63793a",
         837 => x"20000000",
         838 => x"3f0a0000",
         839 => x"3e200000",
         840 => x"68000000",
         841 => x"48656c70",
         842 => x"3a0d0a20",
         843 => x"68202020",
         844 => x"20202020",
         845 => x"20202020",
         846 => x"20202020",
         847 => x"202d2074",
         848 => x"68697320",
         849 => x"68656c70",
         850 => x"0d0a2072",
         851 => x"20202020",
         852 => x"20202020",
         853 => x"20202020",
         854 => x"20202020",
         855 => x"2d207275",
         856 => x"6e206170",
         857 => x"706c6963",
         858 => x"6174696f",
         859 => x"6e0d0a20",
         860 => x"7277203c",
         861 => x"61646472",
         862 => x"3e202020",
         863 => x"20202020",
         864 => x"202d2072",
         865 => x"65616420",
         866 => x"776f7264",
         867 => x"2066726f",
         868 => x"6d206164",
         869 => x"64720d0a",
         870 => x"20777720",
         871 => x"3c616464",
         872 => x"723e203c",
         873 => x"64617461",
         874 => x"3e202d20",
         875 => x"77726974",
         876 => x"6520776f",
         877 => x"72642064",
         878 => x"61746120",
         879 => x"61742061",
         880 => x"6464720d",
         881 => x"0a206477",
         882 => x"203c6164",
         883 => x"64723e20",
         884 => x"20202020",
         885 => x"2020202d",
         886 => x"2064756d",
         887 => x"70203136",
         888 => x"20776f72",
         889 => x"64730d0a",
         890 => x"206e2020",
         891 => x"20202020",
         892 => x"20202020",
         893 => x"20202020",
         894 => x"20202d20",
         895 => x"64756d70",
         896 => x"206e6578",
         897 => x"74203136",
         898 => x"20776f72",
         899 => x"64730000",
         900 => x"72000000",
         901 => x"72772000",
         902 => x"3a200000",
         903 => x"4e6f7420",
         904 => x"6f6e2034",
         905 => x"2d627974",
         906 => x"6520626f",
         907 => x"756e6461",
         908 => x"72792100",
         909 => x"77772000",
         910 => x"64772000",
         911 => x"20200000",
         912 => x"3f3f0000"
            );
end package bootrom_image;
