-- srec2vhdl table generator
-- for input file 'testexceptions.srec'
-- date: Tue Oct 17 16:51:35 2023


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"93828208",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"93804187",
           8 => x"9384019c",
           9 => x"6f000001",
          10 => x"23800000",
          11 => x"93870000",
          12 => x"93801700",
          13 => x"e3ea90fe",
          14 => x"b7070020",
          15 => x"93800700",
          16 => x"93844187",
          17 => x"b7170000",
          18 => x"1389c771",
          19 => x"6f004001",
          20 => x"83470900",
          21 => x"2380f000",
          22 => x"93801000",
          23 => x"13091900",
          24 => x"e3e890fe",
          25 => x"ef00505f",
          26 => x"13060000",
          27 => x"b7070020",
          28 => x"93850700",
          29 => x"13055000",
          30 => x"ef008002",
          31 => x"93000500",
          32 => x"13850000",
          33 => x"ef00c066",
          34 => x"130101ff",
          35 => x"23268100",
          36 => x"13040101",
          37 => x"13000000",
          38 => x"6ff0dfff",
          39 => x"13000000",
          40 => x"130101ff",
          41 => x"23261100",
          42 => x"23248100",
          43 => x"13040101",
          44 => x"93050000",
          45 => x"b7c70100",
          46 => x"13850720",
          47 => x"ef00c053",
          48 => x"97020000",
          49 => x"93820209",
          50 => x"73905230",
          51 => x"b7170000",
          52 => x"13858759",
          53 => x"ef000055",
          54 => x"73000000",
          55 => x"73001000",
          56 => x"b7020030",
          57 => x"03830200",
          58 => x"b7020030",
          59 => x"23806200",
          60 => x"b7020020",
          61 => x"93821200",
          62 => x"03930200",
          63 => x"b7020020",
          64 => x"93821200",
          65 => x"23906200",
          66 => x"b7020020",
          67 => x"93821200",
          68 => x"03a30200",
          69 => x"b7020020",
          70 => x"93821200",
          71 => x"23a06200",
          72 => x"00000000",
          73 => x"b7020020",
          74 => x"67800200",
          75 => x"13000000",
          76 => x"93021000",
          77 => x"67800200",
          78 => x"13000000",
          79 => x"b7170000",
          80 => x"1385475b",
          81 => x"ef00004e",
          82 => x"13000000",
          83 => x"6ff0dfff",
          84 => x"130101fa",
          85 => x"232e1104",
          86 => x"232c5104",
          87 => x"232a6104",
          88 => x"23287104",
          89 => x"23268104",
          90 => x"23249104",
          91 => x"2322a104",
          92 => x"2320b104",
          93 => x"232ec102",
          94 => x"232cd102",
          95 => x"232ae102",
          96 => x"2328f102",
          97 => x"23260103",
          98 => x"23241103",
          99 => x"23222103",
         100 => x"23203103",
         101 => x"232ec101",
         102 => x"232cd101",
         103 => x"232ae101",
         104 => x"2328f101",
         105 => x"13040106",
         106 => x"f3272034",
         107 => x"93800700",
         108 => x"93870000",
         109 => x"13890700",
         110 => x"f3271034",
         111 => x"93800700",
         112 => x"93870000",
         113 => x"93840700",
         114 => x"f3273034",
         115 => x"93800700",
         116 => x"93870000",
         117 => x"93890700",
         118 => x"b7170000",
         119 => x"1385c75b",
         120 => x"ef004044",
         121 => x"93058000",
         122 => x"13050900",
         123 => x"ef008047",
         124 => x"b7170000",
         125 => x"1385475d",
         126 => x"ef00c042",
         127 => x"93058000",
         128 => x"13850400",
         129 => x"ef000046",
         130 => x"b7170000",
         131 => x"1385075e",
         132 => x"ef004041",
         133 => x"93058000",
         134 => x"13850900",
         135 => x"ef008044",
         136 => x"b7170000",
         137 => x"1385c75e",
         138 => x"ef00c03f",
         139 => x"9307b000",
         140 => x"63e6270b",
         141 => x"13172900",
         142 => x"b7170000",
         143 => x"9387c76e",
         144 => x"b307f700",
         145 => x"83a70700",
         146 => x"67800700",
         147 => x"b7170000",
         148 => x"1385075f",
         149 => x"ef00003d",
         150 => x"6f004009",
         151 => x"b7170000",
         152 => x"13850761",
         153 => x"ef00003c",
         154 => x"6f004008",
         155 => x"b7170000",
         156 => x"1385c762",
         157 => x"ef00003b",
         158 => x"6f004007",
         159 => x"b7170000",
         160 => x"13850764",
         161 => x"ef00003a",
         162 => x"6f004006",
         163 => x"b7170000",
         164 => x"13854765",
         165 => x"ef000039",
         166 => x"6f004005",
         167 => x"b7170000",
         168 => x"1385c766",
         169 => x"ef000038",
         170 => x"6f004004",
         171 => x"b7170000",
         172 => x"13850768",
         173 => x"ef000037",
         174 => x"6f004003",
         175 => x"b7170000",
         176 => x"1385c769",
         177 => x"ef000036",
         178 => x"6f004002",
         179 => x"b7170000",
         180 => x"1385076b",
         181 => x"ef000035",
         182 => x"6f004001",
         183 => x"b7170000",
         184 => x"1385876d",
         185 => x"ef000034",
         186 => x"13000000",
         187 => x"b7170000",
         188 => x"1385876e",
         189 => x"ef000033",
         190 => x"93071000",
         191 => x"6316f900",
         192 => x"9304c012",
         193 => x"6f004001",
         194 => x"63160900",
         195 => x"93048013",
         196 => x"6f008000",
         197 => x"93844400",
         198 => x"232694fa",
         199 => x"8327c4fa",
         200 => x"73901734",
         201 => x"13000000",
         202 => x"8320c105",
         203 => x"83228105",
         204 => x"03234105",
         205 => x"83230105",
         206 => x"0324c104",
         207 => x"83248104",
         208 => x"03254104",
         209 => x"83250104",
         210 => x"0326c103",
         211 => x"83268103",
         212 => x"03274103",
         213 => x"83270103",
         214 => x"0328c102",
         215 => x"83288102",
         216 => x"03294102",
         217 => x"83290102",
         218 => x"032ec101",
         219 => x"832e8101",
         220 => x"032f4101",
         221 => x"832f0101",
         222 => x"13010106",
         223 => x"73002030",
         224 => x"13030500",
         225 => x"630a0600",
         226 => x"2300b300",
         227 => x"1306f6ff",
         228 => x"13031300",
         229 => x"e31a06fe",
         230 => x"67800000",
         231 => x"6f000000",
         232 => x"13050000",
         233 => x"67800000",
         234 => x"13050000",
         235 => x"67800000",
         236 => x"130101ff",
         237 => x"23202101",
         238 => x"23261100",
         239 => x"13090600",
         240 => x"6356c002",
         241 => x"23248100",
         242 => x"23229100",
         243 => x"13840500",
         244 => x"b384c500",
         245 => x"03450400",
         246 => x"13041400",
         247 => x"eff05ffc",
         248 => x"e39a84fe",
         249 => x"03248100",
         250 => x"83244100",
         251 => x"8320c100",
         252 => x"13050900",
         253 => x"03290100",
         254 => x"13010101",
         255 => x"67800000",
         256 => x"130101ff",
         257 => x"23202101",
         258 => x"23261100",
         259 => x"13090600",
         260 => x"6356c002",
         261 => x"23248100",
         262 => x"23229100",
         263 => x"13840500",
         264 => x"b384c500",
         265 => x"eff05ff8",
         266 => x"13041400",
         267 => x"a30fa4fe",
         268 => x"e39a84fe",
         269 => x"03248100",
         270 => x"83244100",
         271 => x"8320c100",
         272 => x"13050900",
         273 => x"03290100",
         274 => x"13010101",
         275 => x"67800000",
         276 => x"13051000",
         277 => x"67800000",
         278 => x"130101ff",
         279 => x"23261100",
         280 => x"ef10c008",
         281 => x"8320c100",
         282 => x"93076001",
         283 => x"2320f500",
         284 => x"1305f0ff",
         285 => x"13010101",
         286 => x"67800000",
         287 => x"1305f0ff",
         288 => x"67800000",
         289 => x"b7270000",
         290 => x"23a2f500",
         291 => x"13050000",
         292 => x"67800000",
         293 => x"13051000",
         294 => x"67800000",
         295 => x"13050000",
         296 => x"67800000",
         297 => x"130101fe",
         298 => x"2324c100",
         299 => x"2326d100",
         300 => x"2328e100",
         301 => x"232af100",
         302 => x"232c0101",
         303 => x"232e1101",
         304 => x"1305f0ff",
         305 => x"13010102",
         306 => x"67800000",
         307 => x"130101ff",
         308 => x"23261100",
         309 => x"ef108001",
         310 => x"8320c100",
         311 => x"9307a000",
         312 => x"2320f500",
         313 => x"1305f0ff",
         314 => x"13010101",
         315 => x"67800000",
         316 => x"130101ff",
         317 => x"23261100",
         318 => x"ef00507f",
         319 => x"8320c100",
         320 => x"93072000",
         321 => x"2320f500",
         322 => x"1305f0ff",
         323 => x"13010101",
         324 => x"67800000",
         325 => x"b7270000",
         326 => x"23a2f500",
         327 => x"13050000",
         328 => x"67800000",
         329 => x"130101ff",
         330 => x"23261100",
         331 => x"ef00107c",
         332 => x"8320c100",
         333 => x"9307f001",
         334 => x"2320f500",
         335 => x"1305f0ff",
         336 => x"13010101",
         337 => x"67800000",
         338 => x"130101ff",
         339 => x"23261100",
         340 => x"ef00d079",
         341 => x"8320c100",
         342 => x"9307b000",
         343 => x"2320f500",
         344 => x"1305f0ff",
         345 => x"13010101",
         346 => x"67800000",
         347 => x"130101ff",
         348 => x"23261100",
         349 => x"ef009077",
         350 => x"8320c100",
         351 => x"9307c000",
         352 => x"2320f500",
         353 => x"1305f0ff",
         354 => x"13010101",
         355 => x"67800000",
         356 => x"03a74187",
         357 => x"b7870020",
         358 => x"93870700",
         359 => x"93060040",
         360 => x"b387d740",
         361 => x"630c0700",
         362 => x"3305a700",
         363 => x"63e2a702",
         364 => x"23aaa186",
         365 => x"13050700",
         366 => x"67800000",
         367 => x"9386019c",
         368 => x"1387019c",
         369 => x"23aad186",
         370 => x"3305a700",
         371 => x"e3f2a7fe",
         372 => x"130101ff",
         373 => x"23261100",
         374 => x"ef005071",
         375 => x"8320c100",
         376 => x"9307c000",
         377 => x"2320f500",
         378 => x"1307f0ff",
         379 => x"13050700",
         380 => x"13010101",
         381 => x"67800000",
         382 => x"f32710fc",
         383 => x"63960700",
         384 => x"b7f7fa02",
         385 => x"93870708",
         386 => x"63060500",
         387 => x"33d5a702",
         388 => x"1305f5ff",
         389 => x"b70700f0",
         390 => x"23a6a702",
         391 => x"23a0b702",
         392 => x"67800000",
         393 => x"630e0502",
         394 => x"130101ff",
         395 => x"23248100",
         396 => x"23261100",
         397 => x"13040500",
         398 => x"03450500",
         399 => x"630a0500",
         400 => x"13041400",
         401 => x"ef00c008",
         402 => x"03450400",
         403 => x"e31a05fe",
         404 => x"8320c100",
         405 => x"03248100",
         406 => x"13010101",
         407 => x"67800000",
         408 => x"67800000",
         409 => x"130101fe",
         410 => x"232e1100",
         411 => x"23220100",
         412 => x"23240100",
         413 => x"23060100",
         414 => x"9387f5ff",
         415 => x"13077000",
         416 => x"6376f700",
         417 => x"93077000",
         418 => x"93058000",
         419 => x"13074100",
         420 => x"b307f700",
         421 => x"b385b740",
         422 => x"13069003",
         423 => x"9376f500",
         424 => x"13870603",
         425 => x"6374e600",
         426 => x"13877605",
         427 => x"2380e700",
         428 => x"9387f7ff",
         429 => x"13554500",
         430 => x"e392f5fe",
         431 => x"13054100",
         432 => x"eff05ff6",
         433 => x"8320c101",
         434 => x"13010102",
         435 => x"67800000",
         436 => x"370700f0",
         437 => x"1375f50f",
         438 => x"13070702",
         439 => x"2324a700",
         440 => x"83274700",
         441 => x"93f70701",
         442 => x"e38c07fe",
         443 => x"67800000",
         444 => x"130101ff",
         445 => x"23248100",
         446 => x"23261100",
         447 => x"93070000",
         448 => x"13040500",
         449 => x"63880700",
         450 => x"93050000",
         451 => x"97000000",
         452 => x"e7000000",
         453 => x"83a78187",
         454 => x"63840700",
         455 => x"e7800700",
         456 => x"13050400",
         457 => x"eff09fc7",
         458 => x"13050000",
         459 => x"67800000",
         460 => x"130101ff",
         461 => x"23248100",
         462 => x"23261100",
         463 => x"13040500",
         464 => x"2316b500",
         465 => x"2317c500",
         466 => x"23200500",
         467 => x"23220500",
         468 => x"23240500",
         469 => x"23220506",
         470 => x"23280500",
         471 => x"232a0500",
         472 => x"232c0500",
         473 => x"13068000",
         474 => x"93050000",
         475 => x"1305c505",
         476 => x"eff01fc1",
         477 => x"b7170000",
         478 => x"9387c7a8",
         479 => x"2322f402",
         480 => x"b7170000",
         481 => x"938747ae",
         482 => x"2324f402",
         483 => x"b7170000",
         484 => x"938787b6",
         485 => x"2326f402",
         486 => x"b7170000",
         487 => x"938707bc",
         488 => x"8320c100",
         489 => x"23208402",
         490 => x"2328f402",
         491 => x"03248100",
         492 => x"13010101",
         493 => x"67800000",
         494 => x"b7150000",
         495 => x"37050020",
         496 => x"13868181",
         497 => x"93854541",
         498 => x"13054502",
         499 => x"6f000021",
         500 => x"83254500",
         501 => x"130101ff",
         502 => x"b7070020",
         503 => x"23248100",
         504 => x"23261100",
         505 => x"93878708",
         506 => x"13040500",
         507 => x"6384f500",
         508 => x"ef005042",
         509 => x"83258400",
         510 => x"9387018f",
         511 => x"6386f500",
         512 => x"13050400",
         513 => x"ef001041",
         514 => x"8325c400",
         515 => x"93878195",
         516 => x"638cf500",
         517 => x"13050400",
         518 => x"03248100",
         519 => x"8320c100",
         520 => x"13010101",
         521 => x"6f00103f",
         522 => x"8320c100",
         523 => x"03248100",
         524 => x"13010101",
         525 => x"67800000",
         526 => x"37050020",
         527 => x"130101ff",
         528 => x"9307807b",
         529 => x"13060000",
         530 => x"93054000",
         531 => x"13058508",
         532 => x"23261100",
         533 => x"23acf186",
         534 => x"eff09fed",
         535 => x"13061000",
         536 => x"93059000",
         537 => x"1385018f",
         538 => x"eff09fec",
         539 => x"8320c100",
         540 => x"13062000",
         541 => x"93052001",
         542 => x"13858195",
         543 => x"13010101",
         544 => x"6ff01feb",
         545 => x"13050000",
         546 => x"67800000",
         547 => x"83a78187",
         548 => x"130101ff",
         549 => x"23202101",
         550 => x"23261100",
         551 => x"23248100",
         552 => x"23229100",
         553 => x"13090500",
         554 => x"63940700",
         555 => x"eff0dff8",
         556 => x"93848181",
         557 => x"03a48400",
         558 => x"83a74400",
         559 => x"9387f7ff",
         560 => x"63d80702",
         561 => x"83a70400",
         562 => x"6390070c",
         563 => x"9305c01a",
         564 => x"13050900",
         565 => x"ef00c079",
         566 => x"13040500",
         567 => x"63140508",
         568 => x"23a00400",
         569 => x"9307c000",
         570 => x"2320f900",
         571 => x"6f004005",
         572 => x"0317c400",
         573 => x"63140706",
         574 => x"b707ffff",
         575 => x"93871700",
         576 => x"23220406",
         577 => x"23200400",
         578 => x"23220400",
         579 => x"23240400",
         580 => x"2326f400",
         581 => x"23280400",
         582 => x"232a0400",
         583 => x"232c0400",
         584 => x"13068000",
         585 => x"93050000",
         586 => x"1305c405",
         587 => x"eff05fa5",
         588 => x"232a0402",
         589 => x"232c0402",
         590 => x"23240404",
         591 => x"23260404",
         592 => x"8320c100",
         593 => x"13050400",
         594 => x"03248100",
         595 => x"83244100",
         596 => x"03290100",
         597 => x"13010101",
         598 => x"67800000",
         599 => x"13048406",
         600 => x"6ff0dff5",
         601 => x"93074000",
         602 => x"23200500",
         603 => x"2322f500",
         604 => x"1305c500",
         605 => x"2324a400",
         606 => x"1306001a",
         607 => x"93050000",
         608 => x"eff01fa0",
         609 => x"23a08400",
         610 => x"83a40400",
         611 => x"6ff09ff2",
         612 => x"83270502",
         613 => x"639c0700",
         614 => x"9307007d",
         615 => x"2320f502",
         616 => x"83a78187",
         617 => x"63940700",
         618 => x"6ff01fe9",
         619 => x"67800000",
         620 => x"67800000",
         621 => x"67800000",
         622 => x"13868181",
         623 => x"93058072",
         624 => x"13050000",
         625 => x"6f008001",
         626 => x"b7150000",
         627 => x"13868181",
         628 => x"93854588",
         629 => x"13050000",
         630 => x"6f004000",
         631 => x"130101fd",
         632 => x"23248102",
         633 => x"23202103",
         634 => x"232e3101",
         635 => x"232c4101",
         636 => x"23286101",
         637 => x"23267101",
         638 => x"23261102",
         639 => x"23229102",
         640 => x"232a5101",
         641 => x"93090500",
         642 => x"138a0500",
         643 => x"13040600",
         644 => x"13090000",
         645 => x"130b1000",
         646 => x"930bf0ff",
         647 => x"83248400",
         648 => x"832a4400",
         649 => x"938afaff",
         650 => x"63de0a02",
         651 => x"03240400",
         652 => x"e31604fe",
         653 => x"8320c102",
         654 => x"03248102",
         655 => x"83244102",
         656 => x"8329c101",
         657 => x"032a8101",
         658 => x"832a4101",
         659 => x"032b0101",
         660 => x"832bc100",
         661 => x"13050900",
         662 => x"03290102",
         663 => x"13010103",
         664 => x"67800000",
         665 => x"83d7c400",
         666 => x"637efb00",
         667 => x"8397e400",
         668 => x"638a7701",
         669 => x"93850400",
         670 => x"13850900",
         671 => x"e7000a00",
         672 => x"3369a900",
         673 => x"93848406",
         674 => x"6ff0dff9",
         675 => x"130101ff",
         676 => x"23248100",
         677 => x"13840500",
         678 => x"8395e500",
         679 => x"23261100",
         680 => x"ef008031",
         681 => x"63400502",
         682 => x"83274405",
         683 => x"b387a700",
         684 => x"232af404",
         685 => x"8320c100",
         686 => x"03248100",
         687 => x"13010101",
         688 => x"67800000",
         689 => x"8357c400",
         690 => x"37f7ffff",
         691 => x"1307f7ff",
         692 => x"b3f7e700",
         693 => x"2316f400",
         694 => x"6ff0dffd",
         695 => x"13050000",
         696 => x"67800000",
         697 => x"83d7c500",
         698 => x"130101fe",
         699 => x"232c8100",
         700 => x"232a9100",
         701 => x"23282101",
         702 => x"23263101",
         703 => x"232e1100",
         704 => x"93f70710",
         705 => x"93040500",
         706 => x"13840500",
         707 => x"13090600",
         708 => x"93890600",
         709 => x"638a0700",
         710 => x"8395e500",
         711 => x"93062000",
         712 => x"13060000",
         713 => x"ef004024",
         714 => x"8357c400",
         715 => x"37f7ffff",
         716 => x"1307f7ff",
         717 => x"b3f7e700",
         718 => x"8315e400",
         719 => x"2316f400",
         720 => x"03248101",
         721 => x"8320c101",
         722 => x"93860900",
         723 => x"13060900",
         724 => x"8329c100",
         725 => x"03290101",
         726 => x"13850400",
         727 => x"83244101",
         728 => x"13010102",
         729 => x"6f00402a",
         730 => x"130101ff",
         731 => x"23248100",
         732 => x"13840500",
         733 => x"8395e500",
         734 => x"23261100",
         735 => x"ef00c01e",
         736 => x"1307f0ff",
         737 => x"8357c400",
         738 => x"6312e502",
         739 => x"37f7ffff",
         740 => x"1307f7ff",
         741 => x"b3f7e700",
         742 => x"2316f400",
         743 => x"8320c100",
         744 => x"03248100",
         745 => x"13010101",
         746 => x"67800000",
         747 => x"37170000",
         748 => x"b3e7e700",
         749 => x"2316f400",
         750 => x"232aa404",
         751 => x"6ff01ffe",
         752 => x"8395e500",
         753 => x"6f004000",
         754 => x"130101ff",
         755 => x"23248100",
         756 => x"23229100",
         757 => x"13040500",
         758 => x"13850500",
         759 => x"23261100",
         760 => x"23ae0186",
         761 => x"eff09f89",
         762 => x"9307f0ff",
         763 => x"6318f500",
         764 => x"83a7c187",
         765 => x"63840700",
         766 => x"2320f400",
         767 => x"8320c100",
         768 => x"03248100",
         769 => x"83244100",
         770 => x"13010101",
         771 => x"67800000",
         772 => x"83a70187",
         773 => x"6388a714",
         774 => x"8327c501",
         775 => x"130101fe",
         776 => x"232c8100",
         777 => x"232e1100",
         778 => x"232a9100",
         779 => x"23282101",
         780 => x"23263101",
         781 => x"13040500",
         782 => x"638a0704",
         783 => x"83a7c700",
         784 => x"638c0702",
         785 => x"93040000",
         786 => x"13090008",
         787 => x"8327c401",
         788 => x"83a7c700",
         789 => x"b3879700",
         790 => x"83a50700",
         791 => x"639c050c",
         792 => x"93844400",
         793 => x"e39424ff",
         794 => x"8327c401",
         795 => x"13050400",
         796 => x"83a5c700",
         797 => x"ef000028",
         798 => x"8327c401",
         799 => x"83a50700",
         800 => x"63860500",
         801 => x"13050400",
         802 => x"ef00c026",
         803 => x"83254401",
         804 => x"63860500",
         805 => x"13050400",
         806 => x"ef00c025",
         807 => x"8325c401",
         808 => x"63860500",
         809 => x"13050400",
         810 => x"ef00c024",
         811 => x"83250403",
         812 => x"63860500",
         813 => x"13050400",
         814 => x"ef00c023",
         815 => x"83254403",
         816 => x"63860500",
         817 => x"13050400",
         818 => x"ef00c022",
         819 => x"83258403",
         820 => x"63860500",
         821 => x"13050400",
         822 => x"ef00c021",
         823 => x"83258404",
         824 => x"63860500",
         825 => x"13050400",
         826 => x"ef00c020",
         827 => x"83254404",
         828 => x"63860500",
         829 => x"13050400",
         830 => x"ef00c01f",
         831 => x"8325c402",
         832 => x"63860500",
         833 => x"13050400",
         834 => x"ef00c01e",
         835 => x"83270402",
         836 => x"638c0702",
         837 => x"13050400",
         838 => x"03248101",
         839 => x"8320c101",
         840 => x"83244101",
         841 => x"03290101",
         842 => x"8329c100",
         843 => x"13010102",
         844 => x"67800700",
         845 => x"83a90500",
         846 => x"13050400",
         847 => x"ef00801b",
         848 => x"93850900",
         849 => x"6ff09ff1",
         850 => x"8320c101",
         851 => x"03248101",
         852 => x"83244101",
         853 => x"03290101",
         854 => x"8329c100",
         855 => x"13010102",
         856 => x"67800000",
         857 => x"67800000",
         858 => x"130101ff",
         859 => x"23248100",
         860 => x"23229100",
         861 => x"13040500",
         862 => x"13850500",
         863 => x"93050600",
         864 => x"13860600",
         865 => x"23261100",
         866 => x"23ae0186",
         867 => x"eff00ff1",
         868 => x"9307f0ff",
         869 => x"6318f500",
         870 => x"83a7c187",
         871 => x"63840700",
         872 => x"2320f400",
         873 => x"8320c100",
         874 => x"03248100",
         875 => x"83244100",
         876 => x"13010101",
         877 => x"67800000",
         878 => x"130101ff",
         879 => x"23248100",
         880 => x"23229100",
         881 => x"13040500",
         882 => x"13850500",
         883 => x"93050600",
         884 => x"13860600",
         885 => x"23261100",
         886 => x"23ae0186",
         887 => x"eff04fe2",
         888 => x"9307f0ff",
         889 => x"6318f500",
         890 => x"83a7c187",
         891 => x"63840700",
         892 => x"2320f400",
         893 => x"8320c100",
         894 => x"03248100",
         895 => x"83244100",
         896 => x"13010101",
         897 => x"67800000",
         898 => x"130101ff",
         899 => x"23248100",
         900 => x"23229100",
         901 => x"13040500",
         902 => x"13850500",
         903 => x"93050600",
         904 => x"13860600",
         905 => x"23261100",
         906 => x"23ae0186",
         907 => x"eff04fd8",
         908 => x"9307f0ff",
         909 => x"6318f500",
         910 => x"83a7c187",
         911 => x"63840700",
         912 => x"2320f400",
         913 => x"8320c100",
         914 => x"03248100",
         915 => x"83244100",
         916 => x"13010101",
         917 => x"67800000",
         918 => x"130101ff",
         919 => x"23248100",
         920 => x"23229100",
         921 => x"37140000",
         922 => x"b7140000",
         923 => x"9387c471",
         924 => x"1304c471",
         925 => x"3304f440",
         926 => x"23202101",
         927 => x"23261100",
         928 => x"13542440",
         929 => x"9384c471",
         930 => x"13090000",
         931 => x"63108904",
         932 => x"b7140000",
         933 => x"37140000",
         934 => x"9387c471",
         935 => x"1304c471",
         936 => x"3304f440",
         937 => x"13542440",
         938 => x"9384c471",
         939 => x"13090000",
         940 => x"63188902",
         941 => x"8320c100",
         942 => x"03248100",
         943 => x"83244100",
         944 => x"03290100",
         945 => x"13010101",
         946 => x"67800000",
         947 => x"83a70400",
         948 => x"13091900",
         949 => x"93844400",
         950 => x"e7800700",
         951 => x"6ff01ffb",
         952 => x"83a70400",
         953 => x"13091900",
         954 => x"93844400",
         955 => x"e7800700",
         956 => x"6ff01ffc",
         957 => x"638a050e",
         958 => x"83a7c5ff",
         959 => x"130101fe",
         960 => x"232c8100",
         961 => x"232e1100",
         962 => x"1384c5ff",
         963 => x"63d40700",
         964 => x"3304f400",
         965 => x"2326a100",
         966 => x"ef008031",
         967 => x"83a74188",
         968 => x"0325c100",
         969 => x"639e0700",
         970 => x"23220400",
         971 => x"23a28188",
         972 => x"03248101",
         973 => x"8320c101",
         974 => x"13010102",
         975 => x"6f00802f",
         976 => x"6374f402",
         977 => x"03260400",
         978 => x"b306c400",
         979 => x"639ad700",
         980 => x"83a60700",
         981 => x"83a74700",
         982 => x"b386c600",
         983 => x"2320d400",
         984 => x"2322f400",
         985 => x"6ff09ffc",
         986 => x"13870700",
         987 => x"83a74700",
         988 => x"63840700",
         989 => x"e37af4fe",
         990 => x"83260700",
         991 => x"3306d700",
         992 => x"63188602",
         993 => x"03260400",
         994 => x"b386c600",
         995 => x"2320d700",
         996 => x"3306d700",
         997 => x"e39ec7f8",
         998 => x"03a60700",
         999 => x"83a74700",
        1000 => x"b306d600",
        1001 => x"2320d700",
        1002 => x"2322f700",
        1003 => x"6ff05ff8",
        1004 => x"6378c400",
        1005 => x"9307c000",
        1006 => x"2320f500",
        1007 => x"6ff05ff7",
        1008 => x"03260400",
        1009 => x"b306c400",
        1010 => x"639ad700",
        1011 => x"83a60700",
        1012 => x"83a74700",
        1013 => x"b386c600",
        1014 => x"2320d400",
        1015 => x"2322f400",
        1016 => x"23228700",
        1017 => x"6ff0dff4",
        1018 => x"67800000",
        1019 => x"130101ff",
        1020 => x"23202101",
        1021 => x"83a70188",
        1022 => x"23248100",
        1023 => x"23229100",
        1024 => x"23261100",
        1025 => x"93040500",
        1026 => x"13840500",
        1027 => x"63980700",
        1028 => x"93050000",
        1029 => x"ef000049",
        1030 => x"23a0a188",
        1031 => x"93050400",
        1032 => x"13850400",
        1033 => x"ef000048",
        1034 => x"1309f0ff",
        1035 => x"63122503",
        1036 => x"1304f0ff",
        1037 => x"8320c100",
        1038 => x"13050400",
        1039 => x"03248100",
        1040 => x"83244100",
        1041 => x"03290100",
        1042 => x"13010101",
        1043 => x"67800000",
        1044 => x"13043500",
        1045 => x"1374c4ff",
        1046 => x"e30e85fc",
        1047 => x"b305a440",
        1048 => x"13850400",
        1049 => x"ef000044",
        1050 => x"e31625fd",
        1051 => x"6ff05ffc",
        1052 => x"130101fe",
        1053 => x"232a9100",
        1054 => x"93843500",
        1055 => x"93f4c4ff",
        1056 => x"23282101",
        1057 => x"232e1100",
        1058 => x"232c8100",
        1059 => x"23263101",
        1060 => x"23244101",
        1061 => x"93848400",
        1062 => x"9307c000",
        1063 => x"13090500",
        1064 => x"63f0f40a",
        1065 => x"9304c000",
        1066 => x"63eeb408",
        1067 => x"13050900",
        1068 => x"ef000018",
        1069 => x"83a74188",
        1070 => x"13840700",
        1071 => x"631a040a",
        1072 => x"93850400",
        1073 => x"13050900",
        1074 => x"eff05ff2",
        1075 => x"9307f0ff",
        1076 => x"13040500",
        1077 => x"6316f514",
        1078 => x"03a44188",
        1079 => x"93070400",
        1080 => x"639c0710",
        1081 => x"63040412",
        1082 => x"032a0400",
        1083 => x"93050000",
        1084 => x"13050900",
        1085 => x"330a4401",
        1086 => x"ef00c03a",
        1087 => x"6318aa10",
        1088 => x"83270400",
        1089 => x"13050900",
        1090 => x"b384f440",
        1091 => x"93850400",
        1092 => x"eff0dfed",
        1093 => x"9307f0ff",
        1094 => x"630af50e",
        1095 => x"83270400",
        1096 => x"b3879700",
        1097 => x"2320f400",
        1098 => x"83a74188",
        1099 => x"638e070e",
        1100 => x"03a74700",
        1101 => x"6318870c",
        1102 => x"23a20700",
        1103 => x"6f004006",
        1104 => x"e3d404f6",
        1105 => x"9307c000",
        1106 => x"2320f900",
        1107 => x"13050000",
        1108 => x"8320c101",
        1109 => x"03248101",
        1110 => x"83244101",
        1111 => x"03290101",
        1112 => x"8329c100",
        1113 => x"032a8100",
        1114 => x"13010102",
        1115 => x"67800000",
        1116 => x"83260400",
        1117 => x"b3869640",
        1118 => x"63ca0606",
        1119 => x"1307b000",
        1120 => x"637ad704",
        1121 => x"23209400",
        1122 => x"33079400",
        1123 => x"63908704",
        1124 => x"23a2e188",
        1125 => x"83274400",
        1126 => x"2320d700",
        1127 => x"2322f700",
        1128 => x"13050900",
        1129 => x"ef000009",
        1130 => x"1305b400",
        1131 => x"93074400",
        1132 => x"137585ff",
        1133 => x"3307f540",
        1134 => x"e30cf5f8",
        1135 => x"3304e400",
        1136 => x"b387a740",
        1137 => x"2320f400",
        1138 => x"6ff09ff8",
        1139 => x"23a2e700",
        1140 => x"6ff05ffc",
        1141 => x"03274400",
        1142 => x"63968700",
        1143 => x"23a2e188",
        1144 => x"6ff01ffc",
        1145 => x"23a2e700",
        1146 => x"6ff09ffb",
        1147 => x"93070400",
        1148 => x"03244400",
        1149 => x"6ff09fec",
        1150 => x"13840700",
        1151 => x"83a74700",
        1152 => x"6ff01fee",
        1153 => x"93070700",
        1154 => x"6ff05ff2",
        1155 => x"9307c000",
        1156 => x"2320f900",
        1157 => x"13050900",
        1158 => x"ef00c001",
        1159 => x"6ff01ff3",
        1160 => x"23209500",
        1161 => x"6ff0dff7",
        1162 => x"23220000",
        1163 => x"73001000",
        1164 => x"67800000",
        1165 => x"67800000",
        1166 => x"8397c500",
        1167 => x"130101fe",
        1168 => x"232c8100",
        1169 => x"232a9100",
        1170 => x"232e1100",
        1171 => x"23282101",
        1172 => x"23263101",
        1173 => x"13f78700",
        1174 => x"93040500",
        1175 => x"13840500",
        1176 => x"631a0712",
        1177 => x"03a74500",
        1178 => x"6346e000",
        1179 => x"03a70504",
        1180 => x"6356e010",
        1181 => x"0327c402",
        1182 => x"63020710",
        1183 => x"03a90400",
        1184 => x"93963701",
        1185 => x"23a00400",
        1186 => x"83250402",
        1187 => x"63dc060a",
        1188 => x"03264405",
        1189 => x"8357c400",
        1190 => x"93f74700",
        1191 => x"638e0700",
        1192 => x"83274400",
        1193 => x"3306f640",
        1194 => x"83274403",
        1195 => x"63860700",
        1196 => x"83270404",
        1197 => x"3306f640",
        1198 => x"8327c402",
        1199 => x"83250402",
        1200 => x"93060000",
        1201 => x"13850400",
        1202 => x"e7800700",
        1203 => x"1307f0ff",
        1204 => x"8357c400",
        1205 => x"6312e502",
        1206 => x"83a60400",
        1207 => x"1307d001",
        1208 => x"6362d70a",
        1209 => x"37074020",
        1210 => x"13071700",
        1211 => x"3357d700",
        1212 => x"13771700",
        1213 => x"63080708",
        1214 => x"03270401",
        1215 => x"23220400",
        1216 => x"2320e400",
        1217 => x"13973701",
        1218 => x"635c0700",
        1219 => x"9307f0ff",
        1220 => x"6316f500",
        1221 => x"83a70400",
        1222 => x"63940700",
        1223 => x"232aa404",
        1224 => x"83254403",
        1225 => x"23a02401",
        1226 => x"638a0504",
        1227 => x"93074404",
        1228 => x"6386f500",
        1229 => x"13850400",
        1230 => x"eff0dfbb",
        1231 => x"232a0402",
        1232 => x"6f00c003",
        1233 => x"13060000",
        1234 => x"93061000",
        1235 => x"13850400",
        1236 => x"e7000700",
        1237 => x"9307f0ff",
        1238 => x"13060500",
        1239 => x"e31cf5f2",
        1240 => x"83a70400",
        1241 => x"e38807f2",
        1242 => x"1307d001",
        1243 => x"6386e700",
        1244 => x"13076001",
        1245 => x"6394e706",
        1246 => x"23a02401",
        1247 => x"13050000",
        1248 => x"6f00c006",
        1249 => x"93e70704",
        1250 => x"93970701",
        1251 => x"93d70741",
        1252 => x"6f004005",
        1253 => x"83a90501",
        1254 => x"e38209fe",
        1255 => x"03a90500",
        1256 => x"93f73700",
        1257 => x"23a03501",
        1258 => x"33093941",
        1259 => x"13070000",
        1260 => x"63940700",
        1261 => x"03a74501",
        1262 => x"2324e400",
        1263 => x"e35020fd",
        1264 => x"83278402",
        1265 => x"83250402",
        1266 => x"93060900",
        1267 => x"13860900",
        1268 => x"13850400",
        1269 => x"e7800700",
        1270 => x"6348a002",
        1271 => x"8317c400",
        1272 => x"93e70704",
        1273 => x"2316f400",
        1274 => x"1305f0ff",
        1275 => x"8320c101",
        1276 => x"03248101",
        1277 => x"83244101",
        1278 => x"03290101",
        1279 => x"8329c100",
        1280 => x"13010102",
        1281 => x"67800000",
        1282 => x"b389a900",
        1283 => x"3309a940",
        1284 => x"6ff0dffa",
        1285 => x"83a70501",
        1286 => x"638e0704",
        1287 => x"130101fe",
        1288 => x"232c8100",
        1289 => x"232e1100",
        1290 => x"13040500",
        1291 => x"630c0500",
        1292 => x"83270502",
        1293 => x"63980700",
        1294 => x"2326b100",
        1295 => x"eff04fd5",
        1296 => x"8325c100",
        1297 => x"8397c500",
        1298 => x"638c0700",
        1299 => x"13050400",
        1300 => x"03248101",
        1301 => x"8320c101",
        1302 => x"13010102",
        1303 => x"6ff0dfdd",
        1304 => x"8320c101",
        1305 => x"03248101",
        1306 => x"13050000",
        1307 => x"13010102",
        1308 => x"67800000",
        1309 => x"13050000",
        1310 => x"67800000",
        1311 => x"93050500",
        1312 => x"631e0500",
        1313 => x"b7150000",
        1314 => x"37050020",
        1315 => x"13868181",
        1316 => x"93854541",
        1317 => x"13054502",
        1318 => x"6ff04fd4",
        1319 => x"03a50187",
        1320 => x"6ff05ff7",
        1321 => x"130101ff",
        1322 => x"23248100",
        1323 => x"23229100",
        1324 => x"13040500",
        1325 => x"13850500",
        1326 => x"23261100",
        1327 => x"23ae0186",
        1328 => x"eff00f8d",
        1329 => x"9307f0ff",
        1330 => x"6318f500",
        1331 => x"83a7c187",
        1332 => x"63840700",
        1333 => x"2320f400",
        1334 => x"8320c100",
        1335 => x"03248100",
        1336 => x"83244100",
        1337 => x"13010101",
        1338 => x"67800000",
        1339 => x"03a50187",
        1340 => x"67800000",
        1341 => x"74657374",
        1342 => x"65786365",
        1343 => x"7074696f",
        1344 => x"6e730000",
        1345 => x"54485541",
        1346 => x"53205249",
        1347 => x"53432d56",
        1348 => x"20525633",
        1349 => x"32494d20",
        1350 => x"62617265",
        1351 => x"206d6574",
        1352 => x"616c2070",
        1353 => x"726f6365",
        1354 => x"73736f72",
        1355 => x"00000000",
        1356 => x"54686520",
        1357 => x"48616775",
        1358 => x"6520556e",
        1359 => x"69766572",
        1360 => x"73697479",
        1361 => x"206f6620",
        1362 => x"4170706c",
        1363 => x"69656420",
        1364 => x"53636965",
        1365 => x"6e636573",
        1366 => x"00000000",
        1367 => x"44657061",
        1368 => x"72746d65",
        1369 => x"6e74206f",
        1370 => x"6620456c",
        1371 => x"65637472",
        1372 => x"6963616c",
        1373 => x"20456e67",
        1374 => x"696e6565",
        1375 => x"72696e67",
        1376 => x"00000000",
        1377 => x"4a2e452e",
        1378 => x"4a2e206f",
        1379 => x"70206465",
        1380 => x"6e204272",
        1381 => x"6f757700",
        1382 => x"0d0a4578",
        1383 => x"63657074",
        1384 => x"696f6e20",
        1385 => x"74657374",
        1386 => x"2070726f",
        1387 => x"6772616d",
        1388 => x"0d0a0000",
        1389 => x"446f6e65",
        1390 => x"0d0a0000",
        1391 => x"20457863",
        1392 => x"65707469",
        1393 => x"6f6e2d2d",
        1394 => x"3e206d63",
        1395 => x"61757365",
        1396 => x"3a200000",
        1397 => x"2c206d65",
        1398 => x"70633a20",
        1399 => x"00000000",
        1400 => x"2c206d74",
        1401 => x"76616c3a",
        1402 => x"20000000",
        1403 => x"2c200000",
        1404 => x"496e7374",
        1405 => x"72756374",
        1406 => x"696f6e20",
        1407 => x"61646472",
        1408 => x"65737320",
        1409 => x"6d697361",
        1410 => x"6c69676e",
        1411 => x"65640000",
        1412 => x"496e7374",
        1413 => x"72756374",
        1414 => x"696f6e20",
        1415 => x"61636365",
        1416 => x"73732066",
        1417 => x"61756c74",
        1418 => x"00000000",
        1419 => x"496c6c65",
        1420 => x"67616c20",
        1421 => x"696e7374",
        1422 => x"72756374",
        1423 => x"696f6e00",
        1424 => x"42726561",
        1425 => x"6b706f69",
        1426 => x"6e742028",
        1427 => x"65627265",
        1428 => x"616b2900",
        1429 => x"4c6f6164",
        1430 => x"20616464",
        1431 => x"72657373",
        1432 => x"206d6973",
        1433 => x"616c6967",
        1434 => x"6e656400",
        1435 => x"4c6f6164",
        1436 => x"20616363",
        1437 => x"65737320",
        1438 => x"6661756c",
        1439 => x"74000000",
        1440 => x"53746f72",
        1441 => x"65206164",
        1442 => x"64726573",
        1443 => x"73206d69",
        1444 => x"73616c69",
        1445 => x"676e6564",
        1446 => x"00000000",
        1447 => x"53746f72",
        1448 => x"65206163",
        1449 => x"63657373",
        1450 => x"20666175",
        1451 => x"6c740000",
        1452 => x"456e7669",
        1453 => x"726f6e6d",
        1454 => x"656e7420",
        1455 => x"63616c6c",
        1456 => x"2066726f",
        1457 => x"6d204d2d",
        1458 => x"6d6f6465",
        1459 => x"20286563",
        1460 => x"616c6c29",
        1461 => x"00000000",
        1462 => x"4e6f2064",
        1463 => x"65736372",
        1464 => x"69707469",
        1465 => x"6f6e0000",
        1466 => x"0d0a0000",
        1467 => x"4c020000",
        1468 => x"5c020000",
        1469 => x"6c020000",
        1470 => x"7c020000",
        1471 => x"8c020000",
        1472 => x"9c020000",
        1473 => x"ac020000",
        1474 => x"bc020000",
        1475 => x"dc020000",
        1476 => x"dc020000",
        1477 => x"dc020000",
        1478 => x"cc020000",
        1479 => x"f4140000",
        1480 => x"04150000",
        1481 => x"30150000",
        1482 => x"5c150000",
        1483 => x"84150000",
        1484 => x"00000000",
        1485 => x"00000000",
        1486 => x"03000000",
        1487 => x"88000020",
        1488 => x"00000000",
        1489 => x"88000020",
        1490 => x"f0000020",
        1491 => x"58010020",
        1492 => x"00000000",
        1493 => x"00000000",
        1494 => x"00000000",
        1495 => x"00000000",
        1496 => x"00000000",
        1497 => x"00000000",
        1498 => x"00000000",
        1499 => x"00000000",
        1500 => x"00000000",
        1501 => x"00000000",
        1502 => x"00000000",
        1503 => x"00000000",
        1504 => x"00000000",
        1505 => x"00000000",
        1506 => x"00000000",
        1507 => x"24000020"
            );
end package rom_image;
