-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Thu Jun  5 16:06:25 2025


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382022f",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"37060020",
           9 => x"13050500",
          10 => x"13064607",
          11 => x"637ac500",
          12 => x"b7450000",
          13 => x"3306a640",
          14 => x"938585bb",
          15 => x"ef10c039",
          16 => x"37060020",
          17 => x"13854187",
          18 => x"1306061c",
          19 => x"6378c500",
          20 => x"3306a640",
          21 => x"93050000",
          22 => x"ef104036",
          23 => x"ef20c00d",
          24 => x"b7050020",
          25 => x"93850500",
          26 => x"13060000",
          27 => x"13055000",
          28 => x"ef108047",
          29 => x"ef105005",
          30 => x"6f10003c",
          31 => x"130101fe",
          32 => x"232e1100",
          33 => x"2326a100",
          34 => x"ef100040",
          35 => x"8320c101",
          36 => x"0325c100",
          37 => x"13010102",
          38 => x"67800000",
          39 => x"130101fd",
          40 => x"b7470000",
          41 => x"232c4101",
          42 => x"130a0500",
          43 => x"1385c79c",
          44 => x"23248102",
          45 => x"23229102",
          46 => x"23202103",
          47 => x"232e3101",
          48 => x"83244a08",
          49 => x"23261102",
          50 => x"37390000",
          51 => x"ef10c03d",
          52 => x"13044100",
          53 => x"93070400",
          54 => x"9309c1ff",
          55 => x"13090978",
          56 => x"13f7f400",
          57 => x"3307e900",
          58 => x"03470700",
          59 => x"9387f7ff",
          60 => x"93d44400",
          61 => x"2384e700",
          62 => x"e39437ff",
          63 => x"13054100",
          64 => x"23060100",
          65 => x"ef10403a",
          66 => x"37450000",
          67 => x"1305059e",
          68 => x"ef108039",
          69 => x"03278a08",
          70 => x"9377f700",
          71 => x"b307f900",
          72 => x"83c70700",
          73 => x"1304f4ff",
          74 => x"13574700",
          75 => x"2304f400",
          76 => x"e31434ff",
          77 => x"13054100",
          78 => x"ef100037",
          79 => x"37450000",
          80 => x"1305c59e",
          81 => x"ef104036",
          82 => x"8320c102",
          83 => x"03248102",
          84 => x"83244102",
          85 => x"03290102",
          86 => x"8329c101",
          87 => x"032a8101",
          88 => x"13010103",
          89 => x"67800000",
          90 => x"b70700f0",
          91 => x"03a74760",
          92 => x"93860700",
          93 => x"1377f7fe",
          94 => x"23a2e760",
          95 => x"83a74700",
          96 => x"93c71700",
          97 => x"23a2f600",
          98 => x"67800000",
          99 => x"370700f0",
         100 => x"83274700",
         101 => x"93e70720",
         102 => x"2322f700",
         103 => x"6f000000",
         104 => x"b71700f0",
         105 => x"b71500f0",
         106 => x"938747a0",
         107 => x"938505a0",
         108 => x"83a60700",
         109 => x"03a60500",
         110 => x"03a70700",
         111 => x"e31ad7fe",
         112 => x"b7870100",
         113 => x"b71600f0",
         114 => x"1305f0ff",
         115 => x"9387076a",
         116 => x"23a6a6a0",
         117 => x"b307f600",
         118 => x"23a4a6a0",
         119 => x"33b6c700",
         120 => x"23a4f6a0",
         121 => x"3306e600",
         122 => x"23a6c6a0",
         123 => x"370700f0",
         124 => x"83274700",
         125 => x"93c72700",
         126 => x"2322f700",
         127 => x"67800000",
         128 => x"b70700f0",
         129 => x"03a74710",
         130 => x"b70600f0",
         131 => x"93870710",
         132 => x"13778700",
         133 => x"630a0700",
         134 => x"03a74600",
         135 => x"13478700",
         136 => x"23a2e600",
         137 => x"83a78700",
         138 => x"67800000",
         139 => x"b70700f0",
         140 => x"03a74770",
         141 => x"93860700",
         142 => x"1377f7f0",
         143 => x"23a2e770",
         144 => x"83a74700",
         145 => x"93c74700",
         146 => x"23a2f600",
         147 => x"67800000",
         148 => x"b70700f0",
         149 => x"03a74740",
         150 => x"93860700",
         151 => x"137777ff",
         152 => x"23a2e740",
         153 => x"83a74700",
         154 => x"93c70701",
         155 => x"23a2f600",
         156 => x"67800000",
         157 => x"b70700f0",
         158 => x"03a74720",
         159 => x"93860700",
         160 => x"137777ff",
         161 => x"23a2e720",
         162 => x"83a74700",
         163 => x"93c70702",
         164 => x"23a2f600",
         165 => x"67800000",
         166 => x"b70700f0",
         167 => x"03a74730",
         168 => x"93860700",
         169 => x"137777ff",
         170 => x"23a2e730",
         171 => x"83a74700",
         172 => x"93c70708",
         173 => x"23a2f600",
         174 => x"67800000",
         175 => x"b70700f0",
         176 => x"23ae0700",
         177 => x"03a74700",
         178 => x"13470704",
         179 => x"23a2e700",
         180 => x"67800000",
         181 => x"b71700f0",
         182 => x"23a00790",
         183 => x"370700f0",
         184 => x"83274700",
         185 => x"93c70710",
         186 => x"2322f700",
         187 => x"67800000",
         188 => x"6f000000",
         189 => x"13050000",
         190 => x"67800000",
         191 => x"13050000",
         192 => x"67800000",
         193 => x"130101f7",
         194 => x"23221100",
         195 => x"23242100",
         196 => x"23263100",
         197 => x"23284100",
         198 => x"232a5100",
         199 => x"232c6100",
         200 => x"232e7100",
         201 => x"23208102",
         202 => x"23229102",
         203 => x"2324a102",
         204 => x"2326b102",
         205 => x"2328c102",
         206 => x"232ad102",
         207 => x"232ce102",
         208 => x"232ef102",
         209 => x"23200105",
         210 => x"23221105",
         211 => x"23242105",
         212 => x"23263105",
         213 => x"23284105",
         214 => x"232a5105",
         215 => x"232c6105",
         216 => x"232e7105",
         217 => x"23208107",
         218 => x"23229107",
         219 => x"2324a107",
         220 => x"2326b107",
         221 => x"2328c107",
         222 => x"232ad107",
         223 => x"232ce107",
         224 => x"232ef107",
         225 => x"f3222034",
         226 => x"23205108",
         227 => x"f3221034",
         228 => x"23225108",
         229 => x"83a20200",
         230 => x"23245108",
         231 => x"f3223034",
         232 => x"23265108",
         233 => x"13080100",
         234 => x"ef00400a",
         235 => x"83220108",
         236 => x"63c80200",
         237 => x"73231034",
         238 => x"13034300",
         239 => x"73101334",
         240 => x"1303b000",
         241 => x"63846200",
         242 => x"03258102",
         243 => x"832fc107",
         244 => x"032f8107",
         245 => x"832e4107",
         246 => x"032e0107",
         247 => x"832dc106",
         248 => x"032d8106",
         249 => x"832c4106",
         250 => x"032c0106",
         251 => x"832bc105",
         252 => x"032b8105",
         253 => x"832a4105",
         254 => x"032a0105",
         255 => x"8329c104",
         256 => x"03298104",
         257 => x"83284104",
         258 => x"03280104",
         259 => x"8327c103",
         260 => x"03278103",
         261 => x"83264103",
         262 => x"03260103",
         263 => x"8325c102",
         264 => x"83244102",
         265 => x"03240102",
         266 => x"8323c101",
         267 => x"03238101",
         268 => x"83224101",
         269 => x"03220101",
         270 => x"8321c100",
         271 => x"03218100",
         272 => x"83204100",
         273 => x"13010109",
         274 => x"73002030",
         275 => x"f3272034",
         276 => x"37070080",
         277 => x"1307b701",
         278 => x"6366f720",
         279 => x"130101fe",
         280 => x"37070080",
         281 => x"232e1100",
         282 => x"13072700",
         283 => x"138e0500",
         284 => x"6374f704",
         285 => x"37070080",
         286 => x"1307d7ff",
         287 => x"b387e700",
         288 => x"13078001",
         289 => x"6360f702",
         290 => x"37370000",
         291 => x"93972700",
         292 => x"13074779",
         293 => x"b387e700",
         294 => x"83a70700",
         295 => x"67800700",
         296 => x"eff05fe3",
         297 => x"13060000",
         298 => x"8320c101",
         299 => x"13050600",
         300 => x"13010102",
         301 => x"67800000",
         302 => x"13073000",
         303 => x"6386e704",
         304 => x"1307b000",
         305 => x"e390e7fe",
         306 => x"9307600d",
         307 => x"6380f822",
         308 => x"63e21709",
         309 => x"9307d005",
         310 => x"63ec1719",
         311 => x"93078003",
         312 => x"63f0170b",
         313 => x"938878fc",
         314 => x"93074002",
         315 => x"63ea1709",
         316 => x"b7370000",
         317 => x"9387877f",
         318 => x"93982800",
         319 => x"b388f800",
         320 => x"83a70800",
         321 => x"67800700",
         322 => x"13050800",
         323 => x"eff01fb9",
         324 => x"6ff05ff9",
         325 => x"eff0dfc8",
         326 => x"6ff0dff8",
         327 => x"eff01fda",
         328 => x"6ff05ff8",
         329 => x"eff01fd5",
         330 => x"6ff0dff7",
         331 => x"eff05fd2",
         332 => x"6ff05ff7",
         333 => x"eff05fc3",
         334 => x"6ff0dff6",
         335 => x"eff01fcf",
         336 => x"6ff05ff6",
         337 => x"eff0dfcb",
         338 => x"6ff0dff5",
         339 => x"eff0dfd4",
         340 => x"6ff05ff5",
         341 => x"93073019",
         342 => x"6382f81a",
         343 => x"938808c0",
         344 => x"9307f000",
         345 => x"63ee1701",
         346 => x"b7470000",
         347 => x"9387c788",
         348 => x"93982800",
         349 => x"b388f800",
         350 => x"83a70800",
         351 => x"67800700",
         352 => x"ef10103b",
         353 => x"93078005",
         354 => x"2320f500",
         355 => x"1306f0ff",
         356 => x"6ff09ff1",
         357 => x"b70700f0",
         358 => x"1307f0ff",
         359 => x"23a2e700",
         360 => x"b7270000",
         361 => x"2322fe00",
         362 => x"6ff0dfef",
         363 => x"ef105038",
         364 => x"93079000",
         365 => x"2320f500",
         366 => x"1306f0ff",
         367 => x"6ff0dfee",
         368 => x"ef101037",
         369 => x"9307f001",
         370 => x"2320f500",
         371 => x"1306f0ff",
         372 => x"6ff09fed",
         373 => x"ef10d035",
         374 => x"9307d000",
         375 => x"2320f500",
         376 => x"1306f0ff",
         377 => x"6ff05fec",
         378 => x"ef109034",
         379 => x"93072000",
         380 => x"2320f500",
         381 => x"1306f0ff",
         382 => x"6ff01feb",
         383 => x"e356c0ea",
         384 => x"232c8100",
         385 => x"3384c500",
         386 => x"03450e00",
         387 => x"130e1e00",
         388 => x"2324c100",
         389 => x"2322c101",
         390 => x"eff05fa6",
         391 => x"032e4100",
         392 => x"03268100",
         393 => x"e3128efe",
         394 => x"03248101",
         395 => x"6ff0dfe7",
         396 => x"e35cc0e6",
         397 => x"232c8100",
         398 => x"3384c500",
         399 => x"2324c100",
         400 => x"2322c101",
         401 => x"eff05fa3",
         402 => x"032e4100",
         403 => x"03268100",
         404 => x"2300ae00",
         405 => x"130e1e00",
         406 => x"e3128efe",
         407 => x"03248101",
         408 => x"6ff09fe4",
         409 => x"13060000",
         410 => x"13050600",
         411 => x"67800000",
         412 => x"9307900a",
         413 => x"e396f8f0",
         414 => x"93070000",
         415 => x"2326a100",
         416 => x"13870700",
         417 => x"93860700",
         418 => x"f32710c8",
         419 => x"732710c0",
         420 => x"f32610c8",
         421 => x"e39ad7fe",
         422 => x"37460f00",
         423 => x"13060624",
         424 => x"93060000",
         425 => x"13050700",
         426 => x"93850700",
         427 => x"2324e100",
         428 => x"2322f100",
         429 => x"ef00d00e",
         430 => x"0323c100",
         431 => x"83254100",
         432 => x"37460f00",
         433 => x"2324a300",
         434 => x"03258100",
         435 => x"13060624",
         436 => x"93060000",
         437 => x"23226100",
         438 => x"ef00c04d",
         439 => x"03234100",
         440 => x"2320a300",
         441 => x"2322b300",
         442 => x"6ff0dfdb",
         443 => x"63160508",
         444 => x"37060020",
         445 => x"1306061c",
         446 => x"6ff01fdb",
         447 => x"93070000",
         448 => x"2326b100",
         449 => x"13880700",
         450 => x"13870700",
         451 => x"f32710c8",
         452 => x"732810c0",
         453 => x"732710c8",
         454 => x"e39ae7fe",
         455 => x"37460f00",
         456 => x"13060624",
         457 => x"93060000",
         458 => x"13050800",
         459 => x"93850700",
         460 => x"23240101",
         461 => x"2322f100",
         462 => x"ef009006",
         463 => x"1307803e",
         464 => x"3307e502",
         465 => x"032ec100",
         466 => x"83254100",
         467 => x"03258100",
         468 => x"37460f00",
         469 => x"13060624",
         470 => x"93060000",
         471 => x"2322c101",
         472 => x"2324ee00",
         473 => x"ef000045",
         474 => x"032e4100",
         475 => x"2320ae00",
         476 => x"2322be00",
         477 => x"6ff01fd3",
         478 => x"b7870020",
         479 => x"93870700",
         480 => x"13070040",
         481 => x"b387e740",
         482 => x"6376f500",
         483 => x"13060500",
         484 => x"6ff09fd1",
         485 => x"ef10d019",
         486 => x"9307c000",
         487 => x"2320f500",
         488 => x"1306f0ff",
         489 => x"6ff05fd0",
         490 => x"130e0500",
         491 => x"13830500",
         492 => x"13070000",
         493 => x"63dc0500",
         494 => x"b337a000",
         495 => x"3303b040",
         496 => x"3303f340",
         497 => x"330ea040",
         498 => x"1307f0ff",
         499 => x"63dc0600",
         500 => x"b337c000",
         501 => x"b306d040",
         502 => x"1347f7ff",
         503 => x"b386f640",
         504 => x"3306c040",
         505 => x"13080600",
         506 => x"93850600",
         507 => x"93080e00",
         508 => x"93070300",
         509 => x"63960622",
         510 => x"37450000",
         511 => x"1305c58c",
         512 => x"6374c30e",
         513 => x"b7060100",
         514 => x"6376d60c",
         515 => x"93360610",
         516 => x"93b61600",
         517 => x"93963600",
         518 => x"b35ed600",
         519 => x"3305d501",
         520 => x"03450500",
         521 => x"b306d500",
         522 => x"13050002",
         523 => x"638ea600",
         524 => x"3305d540",
         525 => x"b317a300",
         526 => x"b356de00",
         527 => x"3318a600",
         528 => x"b3e7f600",
         529 => x"b318ae00",
         530 => x"13530801",
         531 => x"33d56702",
         532 => x"13160801",
         533 => x"13560601",
         534 => x"b3f76702",
         535 => x"330ea602",
         536 => x"93960701",
         537 => x"93d70801",
         538 => x"b3e7f600",
         539 => x"63fac701",
         540 => x"b307f800",
         541 => x"63f4c701",
         542 => x"63fa0719",
         543 => x"1305f5ff",
         544 => x"b387c741",
         545 => x"b3d66702",
         546 => x"93980801",
         547 => x"93d80801",
         548 => x"b3f76702",
         549 => x"3306d602",
         550 => x"93970701",
         551 => x"b3e8f800",
         552 => x"63fac800",
         553 => x"b3081801",
         554 => x"63f4c800",
         555 => x"63f60817",
         556 => x"9386f6ff",
         557 => x"13150501",
         558 => x"3365d500",
         559 => x"630a0700",
         560 => x"b337a000",
         561 => x"b305b040",
         562 => x"b385f540",
         563 => x"3305a040",
         564 => x"67800000",
         565 => x"b70e0001",
         566 => x"93068001",
         567 => x"e37ed6f3",
         568 => x"93060001",
         569 => x"6ff05ff3",
         570 => x"93060000",
         571 => x"630c0600",
         572 => x"b7070100",
         573 => x"637af604",
         574 => x"93360610",
         575 => x"93b61600",
         576 => x"93963600",
         577 => x"b357d600",
         578 => x"3305f500",
         579 => x"83470500",
         580 => x"93050002",
         581 => x"b387d700",
         582 => x"6392b704",
         583 => x"b307c340",
         584 => x"93051000",
         585 => x"13530801",
         586 => x"33d56702",
         587 => x"13160801",
         588 => x"13560601",
         589 => x"93d60801",
         590 => x"b3f76702",
         591 => x"330ea602",
         592 => x"93970701",
         593 => x"6ff05ff2",
         594 => x"b7070001",
         595 => x"93068001",
         596 => x"e37af6fa",
         597 => x"93060001",
         598 => x"6ff0dffa",
         599 => x"b385f540",
         600 => x"3318b600",
         601 => x"b356f300",
         602 => x"3313b300",
         603 => x"b357fe00",
         604 => x"b3e76700",
         605 => x"13530801",
         606 => x"b318be00",
         607 => x"b3d56602",
         608 => x"13150801",
         609 => x"13550501",
         610 => x"b3f66602",
         611 => x"330eb502",
         612 => x"13960601",
         613 => x"93d60701",
         614 => x"b3e6c600",
         615 => x"63fac601",
         616 => x"b306d800",
         617 => x"63f4c601",
         618 => x"63f60605",
         619 => x"9385f5ff",
         620 => x"b386c641",
         621 => x"33d66602",
         622 => x"93970701",
         623 => x"93d70701",
         624 => x"b3f66602",
         625 => x"3305c502",
         626 => x"93960601",
         627 => x"b3e7d700",
         628 => x"63faa700",
         629 => x"b307f800",
         630 => x"63f4a700",
         631 => x"63f20703",
         632 => x"1306f6ff",
         633 => x"93950501",
         634 => x"b387a740",
         635 => x"b3e5c500",
         636 => x"6ff05ff3",
         637 => x"9385e5ff",
         638 => x"b3860601",
         639 => x"6ff05ffb",
         640 => x"1306e6ff",
         641 => x"b3870701",
         642 => x"6ff0dffd",
         643 => x"1305e5ff",
         644 => x"b3870701",
         645 => x"6ff0dfe6",
         646 => x"9386e6ff",
         647 => x"6ff09fe9",
         648 => x"6364d318",
         649 => x"b7070100",
         650 => x"63f4f604",
         651 => x"93b50610",
         652 => x"93b51500",
         653 => x"93953500",
         654 => x"b7470000",
         655 => x"33d5b600",
         656 => x"9387c78c",
         657 => x"b387a700",
         658 => x"83c70700",
         659 => x"930e0002",
         660 => x"b387b700",
         661 => x"6398d703",
         662 => x"3335ce00",
         663 => x"13351500",
         664 => x"b3b66600",
         665 => x"3365d500",
         666 => x"93050000",
         667 => x"6ff01fe5",
         668 => x"b7070001",
         669 => x"93058001",
         670 => x"e3f0f6fc",
         671 => x"93050001",
         672 => x"6ff09ffb",
         673 => x"b38efe40",
         674 => x"b355f600",
         675 => x"b396d601",
         676 => x"3358f300",
         677 => x"b3e6d500",
         678 => x"3313d301",
         679 => x"b357fe00",
         680 => x"b3e56700",
         681 => x"13d30601",
         682 => x"b3576802",
         683 => x"13950601",
         684 => x"13550501",
         685 => x"3316d601",
         686 => x"33786802",
         687 => x"330ff502",
         688 => x"93180801",
         689 => x"13d80501",
         690 => x"33681801",
         691 => x"637ae801",
         692 => x"33880601",
         693 => x"6374e801",
         694 => x"637cd80a",
         695 => x"9387f7ff",
         696 => x"3308e841",
         697 => x"b3586802",
         698 => x"93950501",
         699 => x"93d50501",
         700 => x"33786802",
         701 => x"33051503",
         702 => x"13180801",
         703 => x"b3e50501",
         704 => x"63faa500",
         705 => x"b385b600",
         706 => x"63f4a500",
         707 => x"63f8d508",
         708 => x"9388f8ff",
         709 => x"93970701",
         710 => x"13180601",
         711 => x"b385a540",
         712 => x"33e51701",
         713 => x"93980801",
         714 => x"93d80801",
         715 => x"93560501",
         716 => x"13580801",
         717 => x"13560601",
         718 => x"33830803",
         719 => x"33880603",
         720 => x"93570301",
         721 => x"b388c802",
         722 => x"b3880801",
         723 => x"b3871701",
         724 => x"b386c602",
         725 => x"63f60701",
         726 => x"37060100",
         727 => x"b386c600",
         728 => x"13d60701",
         729 => x"b306d600",
         730 => x"63e0d502",
         731 => x"13130301",
         732 => x"93970701",
         733 => x"13530301",
         734 => x"331ede01",
         735 => x"b3876700",
         736 => x"e374feee",
         737 => x"e392d5ee",
         738 => x"1305f5ff",
         739 => x"6ff0dfed",
         740 => x"9387e7ff",
         741 => x"3308d800",
         742 => x"6ff09ff4",
         743 => x"9388e8ff",
         744 => x"b385d500",
         745 => x"6ff01ff7",
         746 => x"93050000",
         747 => x"13050000",
         748 => x"6ff0dfd0",
         749 => x"13070600",
         750 => x"93880600",
         751 => x"13080500",
         752 => x"13830500",
         753 => x"63940624",
         754 => x"b7470000",
         755 => x"9387c78c",
         756 => x"63f4c50e",
         757 => x"b7060100",
         758 => x"6370d60c",
         759 => x"93360610",
         760 => x"93b61600",
         761 => x"93963600",
         762 => x"335ed600",
         763 => x"b387c701",
         764 => x"83c70700",
         765 => x"b387d700",
         766 => x"93060002",
         767 => x"638ed700",
         768 => x"b386f640",
         769 => x"3393d500",
         770 => x"b357f500",
         771 => x"3317d600",
         772 => x"33e36700",
         773 => x"3318d500",
         774 => x"13550701",
         775 => x"b357a302",
         776 => x"93150701",
         777 => x"93d50501",
         778 => x"93560801",
         779 => x"3373a302",
         780 => x"3386f502",
         781 => x"13130301",
         782 => x"b3e66600",
         783 => x"63fac600",
         784 => x"b306d700",
         785 => x"63f4c600",
         786 => x"63f2e606",
         787 => x"9387f7ff",
         788 => x"b386c640",
         789 => x"33d6a602",
         790 => x"13180801",
         791 => x"13580801",
         792 => x"b3f6a602",
         793 => x"b385c502",
         794 => x"93960601",
         795 => x"3368d800",
         796 => x"637ab800",
         797 => x"33080701",
         798 => x"6374b800",
         799 => x"6374e818",
         800 => x"1306f6ff",
         801 => x"93970701",
         802 => x"b3e7c700",
         803 => x"13850700",
         804 => x"93850800",
         805 => x"67800000",
         806 => x"370e0001",
         807 => x"93068001",
         808 => x"e374c6f5",
         809 => x"93060001",
         810 => x"6ff01ff4",
         811 => x"9387e7ff",
         812 => x"b386e600",
         813 => x"6ff0dff9",
         814 => x"93060000",
         815 => x"630c0600",
         816 => x"b7060100",
         817 => x"6378d606",
         818 => x"93360610",
         819 => x"93b61600",
         820 => x"93963600",
         821 => x"b358d600",
         822 => x"b3871701",
         823 => x"83c70700",
         824 => x"b387d700",
         825 => x"93060002",
         826 => x"6390d706",
         827 => x"3386c540",
         828 => x"93081000",
         829 => x"13550701",
         830 => x"b357a602",
         831 => x"93150701",
         832 => x"93d50501",
         833 => x"93560801",
         834 => x"3376a602",
         835 => x"3383f502",
         836 => x"13160601",
         837 => x"b3e6c600",
         838 => x"63fa6600",
         839 => x"b306d700",
         840 => x"63f46600",
         841 => x"63fae60c",
         842 => x"9387f7ff",
         843 => x"b3866640",
         844 => x"6ff05ff2",
         845 => x"b7080001",
         846 => x"93068001",
         847 => x"e37c16f9",
         848 => x"93060001",
         849 => x"6ff01ff9",
         850 => x"3388f640",
         851 => x"33170601",
         852 => x"b3d6f500",
         853 => x"b3950501",
         854 => x"b357f500",
         855 => x"33180501",
         856 => x"13550701",
         857 => x"b3d8a602",
         858 => x"13160701",
         859 => x"13560601",
         860 => x"b3e7b700",
         861 => x"b3f6a602",
         862 => x"33031603",
         863 => x"93950601",
         864 => x"93d60701",
         865 => x"b3e6b600",
         866 => x"63fa6600",
         867 => x"b306d700",
         868 => x"63f46600",
         869 => x"63f6e604",
         870 => x"9388f8ff",
         871 => x"b3866640",
         872 => x"b3d5a602",
         873 => x"93970701",
         874 => x"93d70701",
         875 => x"b3f6a602",
         876 => x"3306b602",
         877 => x"93960601",
         878 => x"b3e7d700",
         879 => x"63fac700",
         880 => x"b307f700",
         881 => x"63f4c700",
         882 => x"63f2e702",
         883 => x"9385f5ff",
         884 => x"93980801",
         885 => x"3386c740",
         886 => x"b3e8b800",
         887 => x"6ff09ff1",
         888 => x"9388e8ff",
         889 => x"b386e600",
         890 => x"6ff05ffb",
         891 => x"9385e5ff",
         892 => x"b387e700",
         893 => x"6ff0dffd",
         894 => x"9387e7ff",
         895 => x"b386e600",
         896 => x"6ff0dff2",
         897 => x"1306e6ff",
         898 => x"6ff0dfe7",
         899 => x"63e4d518",
         900 => x"b7070100",
         901 => x"63f4f604",
         902 => x"93b70610",
         903 => x"93b71700",
         904 => x"93973700",
         905 => x"37470000",
         906 => x"33d8f600",
         907 => x"1307c78c",
         908 => x"33070701",
         909 => x"03470700",
         910 => x"13080002",
         911 => x"3307f700",
         912 => x"63180703",
         913 => x"b337c500",
         914 => x"93b71700",
         915 => x"b3b6b600",
         916 => x"b3e7d700",
         917 => x"93080000",
         918 => x"6ff05fe3",
         919 => x"37070001",
         920 => x"93078001",
         921 => x"e3f0e6fc",
         922 => x"93070001",
         923 => x"6ff09ffb",
         924 => x"3308e840",
         925 => x"b358e600",
         926 => x"b3960601",
         927 => x"b3e8d800",
         928 => x"13de0801",
         929 => x"b3d6e500",
         930 => x"b3d7c603",
         931 => x"13930801",
         932 => x"13530301",
         933 => x"b3950501",
         934 => x"3357e500",
         935 => x"3367b700",
         936 => x"33160601",
         937 => x"b3f6c603",
         938 => x"b30ef302",
         939 => x"93950601",
         940 => x"93560701",
         941 => x"b3e6b600",
         942 => x"63fad601",
         943 => x"b386d800",
         944 => x"63f4d601",
         945 => x"63fc160b",
         946 => x"9387f7ff",
         947 => x"b386d641",
         948 => x"b3d5c603",
         949 => x"13170701",
         950 => x"13570701",
         951 => x"b3f6c603",
         952 => x"3303b302",
         953 => x"93960601",
         954 => x"3367d700",
         955 => x"637a6700",
         956 => x"3387e800",
         957 => x"63746700",
         958 => x"63781709",
         959 => x"9385f5ff",
         960 => x"93970701",
         961 => x"b3e7b700",
         962 => x"33076740",
         963 => x"93950501",
         964 => x"13130601",
         965 => x"93d50501",
         966 => x"93d80701",
         967 => x"13530301",
         968 => x"13560601",
         969 => x"338e6502",
         970 => x"33836802",
         971 => x"93560e01",
         972 => x"b385c502",
         973 => x"b3856500",
         974 => x"b386b600",
         975 => x"b388c802",
         976 => x"63f66600",
         977 => x"37060100",
         978 => x"b388c800",
         979 => x"13d60601",
         980 => x"33061601",
         981 => x"6360c702",
         982 => x"131e0e01",
         983 => x"93960601",
         984 => x"135e0e01",
         985 => x"33150501",
         986 => x"b386c601",
         987 => x"e374d5ee",
         988 => x"e312c7ee",
         989 => x"9387f7ff",
         990 => x"6ff0dfed",
         991 => x"9387e7ff",
         992 => x"b3861601",
         993 => x"6ff09ff4",
         994 => x"9385e5ff",
         995 => x"33071701",
         996 => x"6ff01ff7",
         997 => x"93080000",
         998 => x"93070000",
         999 => x"6ff01fcf",
        1000 => x"13080600",
        1001 => x"93070500",
        1002 => x"13870500",
        1003 => x"63940624",
        1004 => x"b7460000",
        1005 => x"9386c68c",
        1006 => x"63f8c50e",
        1007 => x"b7080100",
        1008 => x"637a160d",
        1009 => x"93380610",
        1010 => x"93b81800",
        1011 => x"93983800",
        1012 => x"33531601",
        1013 => x"b3866600",
        1014 => x"83c60600",
        1015 => x"13030002",
        1016 => x"b3861601",
        1017 => x"b308d340",
        1018 => x"638c6600",
        1019 => x"33971501",
        1020 => x"b356d500",
        1021 => x"33181601",
        1022 => x"33e7e600",
        1023 => x"b3171501",
        1024 => x"13550801",
        1025 => x"b356a702",
        1026 => x"13130801",
        1027 => x"13530301",
        1028 => x"3377a702",
        1029 => x"b3866602",
        1030 => x"93150701",
        1031 => x"13d70701",
        1032 => x"3367b700",
        1033 => x"6370d702",
        1034 => x"3307e800",
        1035 => x"b3350701",
        1036 => x"3336d700",
        1037 => x"93b51500",
        1038 => x"3376b600",
        1039 => x"33060603",
        1040 => x"3307e600",
        1041 => x"3307d740",
        1042 => x"b356a702",
        1043 => x"3377a702",
        1044 => x"b3866602",
        1045 => x"13950701",
        1046 => x"13170701",
        1047 => x"13550501",
        1048 => x"3365e500",
        1049 => x"6370d502",
        1050 => x"3305a800",
        1051 => x"33370501",
        1052 => x"b337d500",
        1053 => x"13371700",
        1054 => x"b3f7e700",
        1055 => x"b3870703",
        1056 => x"3385a700",
        1057 => x"3305d540",
        1058 => x"33551501",
        1059 => x"93050000",
        1060 => x"67800000",
        1061 => x"37030001",
        1062 => x"93088001",
        1063 => x"e37a66f2",
        1064 => x"93080001",
        1065 => x"6ff0dff2",
        1066 => x"13070000",
        1067 => x"630c0600",
        1068 => x"37070100",
        1069 => x"6374e608",
        1070 => x"13370610",
        1071 => x"13371700",
        1072 => x"13173700",
        1073 => x"b358e600",
        1074 => x"b3861601",
        1075 => x"83c60600",
        1076 => x"b386e600",
        1077 => x"13070002",
        1078 => x"b308d740",
        1079 => x"639ae606",
        1080 => x"b386c540",
        1081 => x"93550801",
        1082 => x"33d6b602",
        1083 => x"13130801",
        1084 => x"13530301",
        1085 => x"13d70701",
        1086 => x"b3f6b602",
        1087 => x"33066602",
        1088 => x"93960601",
        1089 => x"3367d700",
        1090 => x"6370c702",
        1091 => x"3307e800",
        1092 => x"33350701",
        1093 => x"b336c700",
        1094 => x"13351500",
        1095 => x"b3f6a600",
        1096 => x"b3860603",
        1097 => x"3387e600",
        1098 => x"3307c740",
        1099 => x"b356b702",
        1100 => x"3377b702",
        1101 => x"b3866602",
        1102 => x"6ff0dff1",
        1103 => x"b7080001",
        1104 => x"13078001",
        1105 => x"e37016f9",
        1106 => x"13070001",
        1107 => x"6ff09ff7",
        1108 => x"33181601",
        1109 => x"33d7d500",
        1110 => x"b3171501",
        1111 => x"b3951501",
        1112 => x"b356d500",
        1113 => x"13550801",
        1114 => x"b3e6b600",
        1115 => x"b355a702",
        1116 => x"131e0801",
        1117 => x"135e0e01",
        1118 => x"3377a702",
        1119 => x"b385c503",
        1120 => x"13160701",
        1121 => x"13d70601",
        1122 => x"3367c700",
        1123 => x"6370b702",
        1124 => x"3307e800",
        1125 => x"33330701",
        1126 => x"3336b700",
        1127 => x"13331300",
        1128 => x"33766600",
        1129 => x"33060603",
        1130 => x"3307e600",
        1131 => x"3307b740",
        1132 => x"3356a702",
        1133 => x"93960601",
        1134 => x"93d60601",
        1135 => x"3377a702",
        1136 => x"3306c603",
        1137 => x"13170701",
        1138 => x"b3e6e600",
        1139 => x"63f0c602",
        1140 => x"b306d800",
        1141 => x"b3b50601",
        1142 => x"33b7c600",
        1143 => x"93b51500",
        1144 => x"3377b700",
        1145 => x"33070703",
        1146 => x"b306d700",
        1147 => x"b386c640",
        1148 => x"6ff05fef",
        1149 => x"63e6d51a",
        1150 => x"37080100",
        1151 => x"63fc0605",
        1152 => x"93b80610",
        1153 => x"93b81800",
        1154 => x"93983800",
        1155 => x"37480000",
        1156 => x"33d31601",
        1157 => x"1308c88c",
        1158 => x"33086800",
        1159 => x"03480800",
        1160 => x"33081801",
        1161 => x"93080002",
        1162 => x"63101805",
        1163 => x"6374c500",
        1164 => x"63fcb600",
        1165 => x"3307c540",
        1166 => x"93070700",
        1167 => x"b386d540",
        1168 => x"3337e500",
        1169 => x"3387e640",
        1170 => x"13850700",
        1171 => x"93050700",
        1172 => x"67800000",
        1173 => x"37080001",
        1174 => x"93088001",
        1175 => x"e3f806fb",
        1176 => x"93080001",
        1177 => x"6ff09ffa",
        1178 => x"b3880841",
        1179 => x"b3961601",
        1180 => x"33530601",
        1181 => x"3363d300",
        1182 => x"33d70501",
        1183 => x"935e0301",
        1184 => x"b356d703",
        1185 => x"131e0301",
        1186 => x"135e0e01",
        1187 => x"b3971501",
        1188 => x"b3550501",
        1189 => x"b3e5f500",
        1190 => x"93d70501",
        1191 => x"33161601",
        1192 => x"33151501",
        1193 => x"3377d703",
        1194 => x"330fde02",
        1195 => x"13170701",
        1196 => x"b3e7e700",
        1197 => x"63fae701",
        1198 => x"b307f300",
        1199 => x"63f4e701",
        1200 => x"63f2670e",
        1201 => x"9386f6ff",
        1202 => x"b387e741",
        1203 => x"33d7d703",
        1204 => x"93950501",
        1205 => x"93d50501",
        1206 => x"b3f7d703",
        1207 => x"330eee02",
        1208 => x"93970701",
        1209 => x"b3e5f500",
        1210 => x"63fac501",
        1211 => x"b305b300",
        1212 => x"63f4c501",
        1213 => x"63fe650a",
        1214 => x"1307f7ff",
        1215 => x"93960601",
        1216 => x"b3e6e600",
        1217 => x"b385c541",
        1218 => x"13170701",
        1219 => x"131e0601",
        1220 => x"93570601",
        1221 => x"13570701",
        1222 => x"93d60601",
        1223 => x"135e0e01",
        1224 => x"b30ec703",
        1225 => x"338ec603",
        1226 => x"3307f702",
        1227 => x"b386f602",
        1228 => x"b307c701",
        1229 => x"13d70e01",
        1230 => x"3307f700",
        1231 => x"6376c701",
        1232 => x"b7070100",
        1233 => x"b386f600",
        1234 => x"93570701",
        1235 => x"939e0e01",
        1236 => x"13170701",
        1237 => x"93de0e01",
        1238 => x"b387d700",
        1239 => x"3307d701",
        1240 => x"63e6f500",
        1241 => x"637ee500",
        1242 => x"639cf500",
        1243 => x"3306c740",
        1244 => x"b336c700",
        1245 => x"b3866600",
        1246 => x"13070600",
        1247 => x"b387d740",
        1248 => x"3307e540",
        1249 => x"3335e500",
        1250 => x"b385f540",
        1251 => x"b385a540",
        1252 => x"33980501",
        1253 => x"33571701",
        1254 => x"3365e800",
        1255 => x"b3d51501",
        1256 => x"67800000",
        1257 => x"9386e6ff",
        1258 => x"b3876700",
        1259 => x"6ff0dff1",
        1260 => x"1307e7ff",
        1261 => x"b3856500",
        1262 => x"6ff05ff4",
        1263 => x"13030500",
        1264 => x"630a0600",
        1265 => x"2300b300",
        1266 => x"1306f6ff",
        1267 => x"13031300",
        1268 => x"e31a06fe",
        1269 => x"67800000",
        1270 => x"13030500",
        1271 => x"630e0600",
        1272 => x"83830500",
        1273 => x"23007300",
        1274 => x"1306f6ff",
        1275 => x"13031300",
        1276 => x"93851500",
        1277 => x"e31606fe",
        1278 => x"67800000",
        1279 => x"630c0602",
        1280 => x"13030500",
        1281 => x"93061000",
        1282 => x"636ab500",
        1283 => x"9306f0ff",
        1284 => x"1307f6ff",
        1285 => x"3303e300",
        1286 => x"b385e500",
        1287 => x"83830500",
        1288 => x"23007300",
        1289 => x"1306f6ff",
        1290 => x"3303d300",
        1291 => x"b385d500",
        1292 => x"e31606fe",
        1293 => x"67800000",
        1294 => x"370700f0",
        1295 => x"13070710",
        1296 => x"83274700",
        1297 => x"93f78700",
        1298 => x"e38c07fe",
        1299 => x"03258700",
        1300 => x"1375f50f",
        1301 => x"67800000",
        1302 => x"f32710fc",
        1303 => x"63960700",
        1304 => x"b7f7fa02",
        1305 => x"93870708",
        1306 => x"63060500",
        1307 => x"33d5a702",
        1308 => x"1305f5ff",
        1309 => x"b70700f0",
        1310 => x"23a6a710",
        1311 => x"23a0b710",
        1312 => x"23a20710",
        1313 => x"67800000",
        1314 => x"370700f0",
        1315 => x"1375f50f",
        1316 => x"13070710",
        1317 => x"2324a700",
        1318 => x"83274700",
        1319 => x"93f70701",
        1320 => x"e38c07fe",
        1321 => x"67800000",
        1322 => x"630e0502",
        1323 => x"130101ff",
        1324 => x"23248100",
        1325 => x"23261100",
        1326 => x"13040500",
        1327 => x"03450500",
        1328 => x"630a0500",
        1329 => x"13041400",
        1330 => x"eff01ffc",
        1331 => x"03450400",
        1332 => x"e31a05fe",
        1333 => x"8320c100",
        1334 => x"03248100",
        1335 => x"13010101",
        1336 => x"67800000",
        1337 => x"67800000",
        1338 => x"130101f9",
        1339 => x"23229106",
        1340 => x"23202107",
        1341 => x"23261106",
        1342 => x"23248106",
        1343 => x"232e3105",
        1344 => x"232a5105",
        1345 => x"23286105",
        1346 => x"23267105",
        1347 => x"23248105",
        1348 => x"23229105",
        1349 => x"2320a105",
        1350 => x"13890500",
        1351 => x"93040500",
        1352 => x"f32a00fc",
        1353 => x"b7070008",
        1354 => x"232c0100",
        1355 => x"232e0100",
        1356 => x"23200102",
        1357 => x"23220102",
        1358 => x"23240102",
        1359 => x"23260102",
        1360 => x"23280102",
        1361 => x"232a0102",
        1362 => x"232c0102",
        1363 => x"232e0102",
        1364 => x"b3fafa00",
        1365 => x"732410fc",
        1366 => x"63160400",
        1367 => x"37f4fa02",
        1368 => x"13040408",
        1369 => x"97f2ffff",
        1370 => x"938202da",
        1371 => x"73905230",
        1372 => x"37c50100",
        1373 => x"13050520",
        1374 => x"93059000",
        1375 => x"eff0dfed",
        1376 => x"b717b7d1",
        1377 => x"93879775",
        1378 => x"b337f402",
        1379 => x"93561400",
        1380 => x"37353e05",
        1381 => x"370600f0",
        1382 => x"13576400",
        1383 => x"130535d6",
        1384 => x"9386f6ff",
        1385 => x"2326d660",
        1386 => x"b725d96f",
        1387 => x"938555d8",
        1388 => x"3337a702",
        1389 => x"93d7d700",
        1390 => x"13051001",
        1391 => x"2320a660",
        1392 => x"9387f7ff",
        1393 => x"2328f670",
        1394 => x"93060600",
        1395 => x"37260000",
        1396 => x"1306f670",
        1397 => x"23a6c670",
        1398 => x"b337b402",
        1399 => x"13576700",
        1400 => x"1307f7ff",
        1401 => x"13860600",
        1402 => x"23a0a670",
        1403 => x"93058070",
        1404 => x"13170701",
        1405 => x"23a0b640",
        1406 => x"13678700",
        1407 => x"2320e620",
        1408 => x"93d73701",
        1409 => x"9387f7ff",
        1410 => x"93970701",
        1411 => x"93e7c700",
        1412 => x"2320f630",
        1413 => x"1307a007",
        1414 => x"93860640",
        1415 => x"232ce600",
        1416 => x"f3224030",
        1417 => x"93e20208",
        1418 => x"73904230",
        1419 => x"f3224030",
        1420 => x"93e28200",
        1421 => x"73904230",
        1422 => x"b7220000",
        1423 => x"93828280",
        1424 => x"73900230",
        1425 => x"b7490000",
        1426 => x"1385c99e",
        1427 => x"eff0dfe5",
        1428 => x"63569002",
        1429 => x"1384f4ff",
        1430 => x"9389c99e",
        1431 => x"9304f0ff",
        1432 => x"03250900",
        1433 => x"1304f4ff",
        1434 => x"13094900",
        1435 => x"eff0dfe3",
        1436 => x"13850900",
        1437 => x"eff05fe3",
        1438 => x"e31494fe",
        1439 => x"37450000",
        1440 => x"1305059f",
        1441 => x"eff05fe2",
        1442 => x"63980a22",
        1443 => x"b7040010",
        1444 => x"37f4eeee",
        1445 => x"b7998888",
        1446 => x"9384f4ff",
        1447 => x"93899988",
        1448 => x"1304f4ee",
        1449 => x"374b0000",
        1450 => x"371c0000",
        1451 => x"37f9eeee",
        1452 => x"130c0c2c",
        1453 => x"1309e9ee",
        1454 => x"6f00c000",
        1455 => x"130cfcff",
        1456 => x"63040c1a",
        1457 => x"93050000",
        1458 => x"13058100",
        1459 => x"ef001030",
        1460 => x"e31605fe",
        1461 => x"832c8100",
        1462 => x"8325c100",
        1463 => x"37160000",
        1464 => x"93d7cc01",
        1465 => x"13974500",
        1466 => x"b307f700",
        1467 => x"33f79700",
        1468 => x"b3f79c00",
        1469 => x"b387e700",
        1470 => x"13d78501",
        1471 => x"b387e700",
        1472 => x"13d7f541",
        1473 => x"1375d700",
        1474 => x"b387a700",
        1475 => x"33b83703",
        1476 => x"137727ff",
        1477 => x"130606e1",
        1478 => x"93060000",
        1479 => x"13850c00",
        1480 => x"130cfcff",
        1481 => x"13583800",
        1482 => x"93184800",
        1483 => x"33880841",
        1484 => x"b3870741",
        1485 => x"b387e700",
        1486 => x"13d7f741",
        1487 => x"b387fc40",
        1488 => x"33b8fc00",
        1489 => x"3387e540",
        1490 => x"33070741",
        1491 => x"33078702",
        1492 => x"33882703",
        1493 => x"33070701",
        1494 => x"33b88702",
        1495 => x"b3878702",
        1496 => x"33070701",
        1497 => x"1358f741",
        1498 => x"13783800",
        1499 => x"b307f800",
        1500 => x"33b80701",
        1501 => x"3308e800",
        1502 => x"1317e801",
        1503 => x"93d72700",
        1504 => x"b307f700",
        1505 => x"93582840",
        1506 => x"13d7c701",
        1507 => x"13934800",
        1508 => x"3307e300",
        1509 => x"33739700",
        1510 => x"33f79700",
        1511 => x"33076700",
        1512 => x"1358f841",
        1513 => x"13d38801",
        1514 => x"33076700",
        1515 => x"1373d800",
        1516 => x"33076700",
        1517 => x"33333703",
        1518 => x"137828ff",
        1519 => x"939b4700",
        1520 => x"b38bfb40",
        1521 => x"939b2b00",
        1522 => x"13533300",
        1523 => x"131e4300",
        1524 => x"33036e40",
        1525 => x"33076740",
        1526 => x"33070701",
        1527 => x"1358f741",
        1528 => x"3387e740",
        1529 => x"33880841",
        1530 => x"b3b8e700",
        1531 => x"33081841",
        1532 => x"33032703",
        1533 => x"33088802",
        1534 => x"b3388702",
        1535 => x"33086800",
        1536 => x"33078702",
        1537 => x"33081801",
        1538 => x"9358f841",
        1539 => x"93f83800",
        1540 => x"3387e800",
        1541 => x"b3381701",
        1542 => x"b3880801",
        1543 => x"9398e801",
        1544 => x"13572700",
        1545 => x"3387e800",
        1546 => x"13184700",
        1547 => x"3307e840",
        1548 => x"13172700",
        1549 => x"338de740",
        1550 => x"efe01ff7",
        1551 => x"83260101",
        1552 => x"13070500",
        1553 => x"33887c41",
        1554 => x"93070d00",
        1555 => x"13860c00",
        1556 => x"93058ba5",
        1557 => x"13058101",
        1558 => x"ef008047",
        1559 => x"13058101",
        1560 => x"eff09fc4",
        1561 => x"e3100ce6",
        1562 => x"63940a00",
        1563 => x"73001000",
        1564 => x"b70700f0",
        1565 => x"1307f00f",
        1566 => x"23a4e740",
        1567 => x"370700f0",
        1568 => x"83260720",
        1569 => x"13060009",
        1570 => x"93070700",
        1571 => x"93e60630",
        1572 => x"2320d720",
        1573 => x"2324c720",
        1574 => x"83260730",
        1575 => x"371700f0",
        1576 => x"93e60630",
        1577 => x"23a0d730",
        1578 => x"23a4c730",
        1579 => x"93071000",
        1580 => x"2320f790",
        1581 => x"6ff05fdf",
        1582 => x"37450000",
        1583 => x"130505a2",
        1584 => x"eff09fbe",
        1585 => x"6ff09fdc",
        1586 => x"130101ff",
        1587 => x"23248100",
        1588 => x"23261100",
        1589 => x"93070000",
        1590 => x"13040500",
        1591 => x"63880700",
        1592 => x"93050000",
        1593 => x"97000000",
        1594 => x"e7000000",
        1595 => x"83a74187",
        1596 => x"63840700",
        1597 => x"e7800700",
        1598 => x"13050400",
        1599 => x"ef101044",
        1600 => x"13050000",
        1601 => x"67800000",
        1602 => x"130101ff",
        1603 => x"23248100",
        1604 => x"23261100",
        1605 => x"13040500",
        1606 => x"2316b500",
        1607 => x"2317c500",
        1608 => x"23200500",
        1609 => x"23220500",
        1610 => x"23240500",
        1611 => x"23220506",
        1612 => x"23280500",
        1613 => x"232a0500",
        1614 => x"232c0500",
        1615 => x"13068000",
        1616 => x"93050000",
        1617 => x"1305c505",
        1618 => x"eff05fa7",
        1619 => x"b7270000",
        1620 => x"938747d4",
        1621 => x"2322f402",
        1622 => x"b7270000",
        1623 => x"9387c7d9",
        1624 => x"2324f402",
        1625 => x"b7270000",
        1626 => x"938707e2",
        1627 => x"2326f402",
        1628 => x"b7270000",
        1629 => x"938787e7",
        1630 => x"8320c100",
        1631 => x"23208402",
        1632 => x"2328f402",
        1633 => x"03248100",
        1634 => x"13010101",
        1635 => x"67800000",
        1636 => x"b7350000",
        1637 => x"37050020",
        1638 => x"13868181",
        1639 => x"9385c52d",
        1640 => x"13054502",
        1641 => x"6f00c021",
        1642 => x"83254500",
        1643 => x"130101ff",
        1644 => x"b7070020",
        1645 => x"23248100",
        1646 => x"23261100",
        1647 => x"93878708",
        1648 => x"13040500",
        1649 => x"6384f500",
        1650 => x"ef105011",
        1651 => x"83258400",
        1652 => x"9387018f",
        1653 => x"6386f500",
        1654 => x"13050400",
        1655 => x"ef101010",
        1656 => x"8325c400",
        1657 => x"93878195",
        1658 => x"638cf500",
        1659 => x"13050400",
        1660 => x"03248100",
        1661 => x"8320c100",
        1662 => x"13010101",
        1663 => x"6f10100e",
        1664 => x"8320c100",
        1665 => x"03248100",
        1666 => x"13010101",
        1667 => x"67800000",
        1668 => x"b7270000",
        1669 => x"37050020",
        1670 => x"130101ff",
        1671 => x"93870799",
        1672 => x"13060000",
        1673 => x"93054000",
        1674 => x"13058508",
        1675 => x"23261100",
        1676 => x"23aaf186",
        1677 => x"eff05fed",
        1678 => x"13061000",
        1679 => x"93059000",
        1680 => x"1385018f",
        1681 => x"eff05fec",
        1682 => x"8320c100",
        1683 => x"13062000",
        1684 => x"93052001",
        1685 => x"13858195",
        1686 => x"13010101",
        1687 => x"6ff0dfea",
        1688 => x"13050000",
        1689 => x"67800000",
        1690 => x"83a74187",
        1691 => x"130101ff",
        1692 => x"23202101",
        1693 => x"23261100",
        1694 => x"23248100",
        1695 => x"23229100",
        1696 => x"13090500",
        1697 => x"63940700",
        1698 => x"eff09ff8",
        1699 => x"93848181",
        1700 => x"03a48400",
        1701 => x"83a74400",
        1702 => x"9387f7ff",
        1703 => x"63d80702",
        1704 => x"03a40400",
        1705 => x"6310040c",
        1706 => x"9305c01a",
        1707 => x"13050900",
        1708 => x"ef00900a",
        1709 => x"13040500",
        1710 => x"63140508",
        1711 => x"23a00400",
        1712 => x"9307c000",
        1713 => x"2320f900",
        1714 => x"6f004005",
        1715 => x"0317c400",
        1716 => x"63140706",
        1717 => x"b707ffff",
        1718 => x"93871700",
        1719 => x"23220406",
        1720 => x"23200400",
        1721 => x"23220400",
        1722 => x"23240400",
        1723 => x"2326f400",
        1724 => x"23280400",
        1725 => x"232a0400",
        1726 => x"232c0400",
        1727 => x"13068000",
        1728 => x"93050000",
        1729 => x"1305c405",
        1730 => x"eff05f8b",
        1731 => x"232a0402",
        1732 => x"232c0402",
        1733 => x"23240404",
        1734 => x"23260404",
        1735 => x"8320c100",
        1736 => x"13050400",
        1737 => x"03248100",
        1738 => x"83244100",
        1739 => x"03290100",
        1740 => x"13010101",
        1741 => x"67800000",
        1742 => x"13048406",
        1743 => x"6ff0dff5",
        1744 => x"93074000",
        1745 => x"23200500",
        1746 => x"2322f500",
        1747 => x"1305c500",
        1748 => x"2324a400",
        1749 => x"1306001a",
        1750 => x"93050000",
        1751 => x"eff01f86",
        1752 => x"23a08400",
        1753 => x"93040400",
        1754 => x"6ff09ff2",
        1755 => x"83270502",
        1756 => x"639e0700",
        1757 => x"b7270000",
        1758 => x"9387879a",
        1759 => x"2320f502",
        1760 => x"83a74187",
        1761 => x"63940700",
        1762 => x"6ff09fe8",
        1763 => x"67800000",
        1764 => x"67800000",
        1765 => x"67800000",
        1766 => x"b7250000",
        1767 => x"13868181",
        1768 => x"93850590",
        1769 => x"13050000",
        1770 => x"6f008001",
        1771 => x"b7250000",
        1772 => x"13868181",
        1773 => x"938505a6",
        1774 => x"13050000",
        1775 => x"6f004000",
        1776 => x"130101fd",
        1777 => x"23248102",
        1778 => x"23202103",
        1779 => x"232e3101",
        1780 => x"232c4101",
        1781 => x"232a5101",
        1782 => x"23261102",
        1783 => x"23229102",
        1784 => x"130a0500",
        1785 => x"938a0500",
        1786 => x"13040000",
        1787 => x"13091000",
        1788 => x"9309f0ff",
        1789 => x"83258600",
        1790 => x"83244600",
        1791 => x"9384f4ff",
        1792 => x"63da0402",
        1793 => x"03260600",
        1794 => x"e31606fe",
        1795 => x"8320c102",
        1796 => x"13050400",
        1797 => x"03248102",
        1798 => x"83244102",
        1799 => x"03290102",
        1800 => x"8329c101",
        1801 => x"032a8101",
        1802 => x"832a4101",
        1803 => x"13010103",
        1804 => x"67800000",
        1805 => x"83d7c500",
        1806 => x"6374f902",
        1807 => x"8397e500",
        1808 => x"63803703",
        1809 => x"13050a00",
        1810 => x"2326c100",
        1811 => x"2324b100",
        1812 => x"e7800a00",
        1813 => x"0326c100",
        1814 => x"83258100",
        1815 => x"3364a400",
        1816 => x"93858506",
        1817 => x"6ff09ff9",
        1818 => x"130101f6",
        1819 => x"232af108",
        1820 => x"b7070080",
        1821 => x"9387f7ff",
        1822 => x"232ef100",
        1823 => x"2328f100",
        1824 => x"b707ffff",
        1825 => x"2326d108",
        1826 => x"2324b100",
        1827 => x"232cb100",
        1828 => x"93878720",
        1829 => x"9306c108",
        1830 => x"93058100",
        1831 => x"232e1106",
        1832 => x"232af100",
        1833 => x"2328e108",
        1834 => x"232c0109",
        1835 => x"232e1109",
        1836 => x"23260106",
        1837 => x"2322d100",
        1838 => x"ef00103a",
        1839 => x"83278100",
        1840 => x"23800700",
        1841 => x"8320c107",
        1842 => x"1301010a",
        1843 => x"67800000",
        1844 => x"130101f6",
        1845 => x"232af108",
        1846 => x"b7070080",
        1847 => x"9387f7ff",
        1848 => x"232ef100",
        1849 => x"2328f100",
        1850 => x"b707ffff",
        1851 => x"93878720",
        1852 => x"232af100",
        1853 => x"2324a100",
        1854 => x"232ca100",
        1855 => x"03a50187",
        1856 => x"2324c108",
        1857 => x"2326d108",
        1858 => x"13860500",
        1859 => x"93068108",
        1860 => x"93058100",
        1861 => x"232e1106",
        1862 => x"2328e108",
        1863 => x"232c0109",
        1864 => x"232e1109",
        1865 => x"23260106",
        1866 => x"2322d100",
        1867 => x"ef00d032",
        1868 => x"83278100",
        1869 => x"23800700",
        1870 => x"8320c107",
        1871 => x"1301010a",
        1872 => x"67800000",
        1873 => x"130101ff",
        1874 => x"23248100",
        1875 => x"13840500",
        1876 => x"8395e500",
        1877 => x"23261100",
        1878 => x"ef008033",
        1879 => x"63400502",
        1880 => x"83274405",
        1881 => x"b387a700",
        1882 => x"232af404",
        1883 => x"8320c100",
        1884 => x"03248100",
        1885 => x"13010101",
        1886 => x"67800000",
        1887 => x"8357c400",
        1888 => x"37f7ffff",
        1889 => x"1307f7ff",
        1890 => x"b3f7e700",
        1891 => x"2316f400",
        1892 => x"6ff0dffd",
        1893 => x"13050000",
        1894 => x"67800000",
        1895 => x"83d7c500",
        1896 => x"130101fe",
        1897 => x"232c8100",
        1898 => x"232a9100",
        1899 => x"23282101",
        1900 => x"23263101",
        1901 => x"232e1100",
        1902 => x"93f70710",
        1903 => x"93040500",
        1904 => x"13840500",
        1905 => x"13090600",
        1906 => x"93890600",
        1907 => x"638a0700",
        1908 => x"8395e500",
        1909 => x"93062000",
        1910 => x"13060000",
        1911 => x"ef004026",
        1912 => x"8357c400",
        1913 => x"37f7ffff",
        1914 => x"1307f7ff",
        1915 => x"b3f7e700",
        1916 => x"8315e400",
        1917 => x"2316f400",
        1918 => x"03248101",
        1919 => x"8320c101",
        1920 => x"93860900",
        1921 => x"13060900",
        1922 => x"8329c100",
        1923 => x"03290101",
        1924 => x"13850400",
        1925 => x"83244101",
        1926 => x"13010102",
        1927 => x"6f00402c",
        1928 => x"130101ff",
        1929 => x"23248100",
        1930 => x"13840500",
        1931 => x"8395e500",
        1932 => x"23261100",
        1933 => x"ef00c020",
        1934 => x"1307f0ff",
        1935 => x"8317c400",
        1936 => x"6312e502",
        1937 => x"13070580",
        1938 => x"13070780",
        1939 => x"b3f7e700",
        1940 => x"2316f400",
        1941 => x"8320c100",
        1942 => x"03248100",
        1943 => x"13010101",
        1944 => x"67800000",
        1945 => x"37170000",
        1946 => x"b3e7e700",
        1947 => x"2316f400",
        1948 => x"232aa404",
        1949 => x"6ff01ffe",
        1950 => x"8395e500",
        1951 => x"6f004000",
        1952 => x"130101ff",
        1953 => x"23248100",
        1954 => x"23229100",
        1955 => x"93040500",
        1956 => x"13850500",
        1957 => x"23261100",
        1958 => x"23ac0186",
        1959 => x"ef100066",
        1960 => x"9307f0ff",
        1961 => x"6318f500",
        1962 => x"83a78187",
        1963 => x"63840700",
        1964 => x"23a0f400",
        1965 => x"8320c100",
        1966 => x"03248100",
        1967 => x"83244100",
        1968 => x"13010101",
        1969 => x"67800000",
        1970 => x"83a70187",
        1971 => x"6388a716",
        1972 => x"8327c501",
        1973 => x"130101fe",
        1974 => x"232c8100",
        1975 => x"232e1100",
        1976 => x"232a9100",
        1977 => x"23282101",
        1978 => x"23263101",
        1979 => x"13040500",
        1980 => x"63840708",
        1981 => x"83a7c700",
        1982 => x"638c0702",
        1983 => x"93040000",
        1984 => x"13090008",
        1985 => x"8327c401",
        1986 => x"83a7c700",
        1987 => x"b3879700",
        1988 => x"83a50700",
        1989 => x"63980504",
        1990 => x"93844400",
        1991 => x"e39424ff",
        1992 => x"8327c401",
        1993 => x"13050400",
        1994 => x"83a5c700",
        1995 => x"ef00002b",
        1996 => x"8327c401",
        1997 => x"83a50700",
        1998 => x"63860500",
        1999 => x"13050400",
        2000 => x"ef00c029",
        2001 => x"8327c401",
        2002 => x"83a48700",
        2003 => x"63860402",
        2004 => x"93850400",
        2005 => x"13050400",
        2006 => x"83a40400",
        2007 => x"ef000028",
        2008 => x"6ff0dffe",
        2009 => x"83a90500",
        2010 => x"13050400",
        2011 => x"ef000027",
        2012 => x"93850900",
        2013 => x"6ff01ffa",
        2014 => x"83254401",
        2015 => x"63860500",
        2016 => x"13050400",
        2017 => x"ef008025",
        2018 => x"8325c401",
        2019 => x"63860500",
        2020 => x"13050400",
        2021 => x"ef008024",
        2022 => x"83250403",
        2023 => x"63860500",
        2024 => x"13050400",
        2025 => x"ef008023",
        2026 => x"83254403",
        2027 => x"63860500",
        2028 => x"13050400",
        2029 => x"ef008022",
        2030 => x"83258403",
        2031 => x"63860500",
        2032 => x"13050400",
        2033 => x"ef008021",
        2034 => x"83258404",
        2035 => x"63860500",
        2036 => x"13050400",
        2037 => x"ef008020",
        2038 => x"83254404",
        2039 => x"63860500",
        2040 => x"13050400",
        2041 => x"ef00801f",
        2042 => x"8325c402",
        2043 => x"63860500",
        2044 => x"13050400",
        2045 => x"ef00801e",
        2046 => x"83270402",
        2047 => x"63820702",
        2048 => x"13050400",
        2049 => x"03248101",
        2050 => x"8320c101",
        2051 => x"83244101",
        2052 => x"03290101",
        2053 => x"8329c100",
        2054 => x"13010102",
        2055 => x"67800700",
        2056 => x"8320c101",
        2057 => x"03248101",
        2058 => x"83244101",
        2059 => x"03290101",
        2060 => x"8329c100",
        2061 => x"13010102",
        2062 => x"67800000",
        2063 => x"67800000",
        2064 => x"130101ff",
        2065 => x"23248100",
        2066 => x"23229100",
        2067 => x"93040500",
        2068 => x"13850500",
        2069 => x"93050600",
        2070 => x"13860600",
        2071 => x"23261100",
        2072 => x"23ac0186",
        2073 => x"ef10c057",
        2074 => x"9307f0ff",
        2075 => x"6318f500",
        2076 => x"83a78187",
        2077 => x"63840700",
        2078 => x"23a0f400",
        2079 => x"8320c100",
        2080 => x"03248100",
        2081 => x"83244100",
        2082 => x"13010101",
        2083 => x"67800000",
        2084 => x"130101ff",
        2085 => x"23248100",
        2086 => x"23229100",
        2087 => x"93040500",
        2088 => x"13850500",
        2089 => x"93050600",
        2090 => x"13860600",
        2091 => x"23261100",
        2092 => x"23ac0186",
        2093 => x"ef10c056",
        2094 => x"9307f0ff",
        2095 => x"6318f500",
        2096 => x"83a78187",
        2097 => x"63840700",
        2098 => x"23a0f400",
        2099 => x"8320c100",
        2100 => x"03248100",
        2101 => x"83244100",
        2102 => x"13010101",
        2103 => x"67800000",
        2104 => x"130101ff",
        2105 => x"23248100",
        2106 => x"23229100",
        2107 => x"93040500",
        2108 => x"13850500",
        2109 => x"93050600",
        2110 => x"13860600",
        2111 => x"23261100",
        2112 => x"23ac0186",
        2113 => x"ef10405c",
        2114 => x"9307f0ff",
        2115 => x"6318f500",
        2116 => x"83a78187",
        2117 => x"63840700",
        2118 => x"23a0f400",
        2119 => x"8320c100",
        2120 => x"03248100",
        2121 => x"83244100",
        2122 => x"13010101",
        2123 => x"67800000",
        2124 => x"03a50187",
        2125 => x"67800000",
        2126 => x"130101ff",
        2127 => x"23248100",
        2128 => x"23229100",
        2129 => x"37440000",
        2130 => x"b7440000",
        2131 => x"130484bb",
        2132 => x"938484bb",
        2133 => x"b3848440",
        2134 => x"23202101",
        2135 => x"23261100",
        2136 => x"93d42440",
        2137 => x"13090000",
        2138 => x"631e9902",
        2139 => x"37440000",
        2140 => x"b7440000",
        2141 => x"130484bb",
        2142 => x"938484bb",
        2143 => x"b3848440",
        2144 => x"93d42440",
        2145 => x"13090000",
        2146 => x"63189902",
        2147 => x"8320c100",
        2148 => x"03248100",
        2149 => x"83244100",
        2150 => x"03290100",
        2151 => x"13010101",
        2152 => x"67800000",
        2153 => x"83270400",
        2154 => x"13091900",
        2155 => x"13044400",
        2156 => x"e7800700",
        2157 => x"6ff05ffb",
        2158 => x"83270400",
        2159 => x"13091900",
        2160 => x"13044400",
        2161 => x"e7800700",
        2162 => x"6ff01ffc",
        2163 => x"13860500",
        2164 => x"93050500",
        2165 => x"03a50187",
        2166 => x"6f10801b",
        2167 => x"638a050e",
        2168 => x"83a7c5ff",
        2169 => x"130101fe",
        2170 => x"232c8100",
        2171 => x"232e1100",
        2172 => x"1384c5ff",
        2173 => x"63d40700",
        2174 => x"3304f400",
        2175 => x"2326a100",
        2176 => x"ef004031",
        2177 => x"83a70188",
        2178 => x"0325c100",
        2179 => x"639e0700",
        2180 => x"23220400",
        2181 => x"23a08188",
        2182 => x"03248101",
        2183 => x"8320c101",
        2184 => x"13010102",
        2185 => x"6f00402f",
        2186 => x"6374f402",
        2187 => x"03260400",
        2188 => x"b306c400",
        2189 => x"639ad700",
        2190 => x"83a60700",
        2191 => x"83a74700",
        2192 => x"b386c600",
        2193 => x"2320d400",
        2194 => x"2322f400",
        2195 => x"6ff09ffc",
        2196 => x"13870700",
        2197 => x"83a74700",
        2198 => x"63840700",
        2199 => x"e37af4fe",
        2200 => x"83260700",
        2201 => x"3306d700",
        2202 => x"63188602",
        2203 => x"03260400",
        2204 => x"b386c600",
        2205 => x"2320d700",
        2206 => x"3306d700",
        2207 => x"e39ec7f8",
        2208 => x"03a60700",
        2209 => x"83a74700",
        2210 => x"b306d600",
        2211 => x"2320d700",
        2212 => x"2322f700",
        2213 => x"6ff05ff8",
        2214 => x"6378c400",
        2215 => x"9307c000",
        2216 => x"2320f500",
        2217 => x"6ff05ff7",
        2218 => x"03260400",
        2219 => x"b306c400",
        2220 => x"639ad700",
        2221 => x"83a60700",
        2222 => x"83a74700",
        2223 => x"b386c600",
        2224 => x"2320d400",
        2225 => x"2322f400",
        2226 => x"23228700",
        2227 => x"6ff0dff4",
        2228 => x"67800000",
        2229 => x"130101ff",
        2230 => x"23248100",
        2231 => x"83a7c187",
        2232 => x"23229100",
        2233 => x"23202101",
        2234 => x"23261100",
        2235 => x"13090500",
        2236 => x"93840500",
        2237 => x"63980700",
        2238 => x"93050000",
        2239 => x"ef10000e",
        2240 => x"23aea186",
        2241 => x"93850400",
        2242 => x"13050900",
        2243 => x"ef10000d",
        2244 => x"9304f0ff",
        2245 => x"63129502",
        2246 => x"1304f0ff",
        2247 => x"8320c100",
        2248 => x"13050400",
        2249 => x"03248100",
        2250 => x"83244100",
        2251 => x"03290100",
        2252 => x"13010101",
        2253 => x"67800000",
        2254 => x"13043500",
        2255 => x"1374c4ff",
        2256 => x"e30e85fc",
        2257 => x"b305a440",
        2258 => x"13050900",
        2259 => x"ef100009",
        2260 => x"e31695fc",
        2261 => x"6ff05ffc",
        2262 => x"130101fe",
        2263 => x"232a9100",
        2264 => x"93843500",
        2265 => x"93f4c4ff",
        2266 => x"232e1100",
        2267 => x"232c8100",
        2268 => x"23282101",
        2269 => x"23263101",
        2270 => x"23244101",
        2271 => x"93848400",
        2272 => x"9307c000",
        2273 => x"63f4f400",
        2274 => x"93840700",
        2275 => x"63c40400",
        2276 => x"63f8b402",
        2277 => x"9307c000",
        2278 => x"2320f500",
        2279 => x"13050000",
        2280 => x"8320c101",
        2281 => x"03248101",
        2282 => x"83244101",
        2283 => x"03290101",
        2284 => x"8329c100",
        2285 => x"032a8100",
        2286 => x"13010102",
        2287 => x"67800000",
        2288 => x"13090500",
        2289 => x"ef000015",
        2290 => x"83a70188",
        2291 => x"13840700",
        2292 => x"63100408",
        2293 => x"93850400",
        2294 => x"13050900",
        2295 => x"eff09fef",
        2296 => x"9307f0ff",
        2297 => x"13040500",
        2298 => x"6312f512",
        2299 => x"03a40188",
        2300 => x"93070400",
        2301 => x"6392070e",
        2302 => x"63000410",
        2303 => x"032a0400",
        2304 => x"93050000",
        2305 => x"13050900",
        2306 => x"330a4401",
        2307 => x"ef00107d",
        2308 => x"6314aa0e",
        2309 => x"83270400",
        2310 => x"13050900",
        2311 => x"b384f440",
        2312 => x"93850400",
        2313 => x"eff01feb",
        2314 => x"9307f0ff",
        2315 => x"6306f50c",
        2316 => x"83270400",
        2317 => x"b3879700",
        2318 => x"2320f400",
        2319 => x"83a70188",
        2320 => x"03a74700",
        2321 => x"6310070a",
        2322 => x"23a00188",
        2323 => x"6f004003",
        2324 => x"83260400",
        2325 => x"b3869640",
        2326 => x"63ca0606",
        2327 => x"1307b000",
        2328 => x"637ad704",
        2329 => x"23209400",
        2330 => x"33079400",
        2331 => x"63908704",
        2332 => x"23a0e188",
        2333 => x"83274400",
        2334 => x"2320d700",
        2335 => x"2322f700",
        2336 => x"13050900",
        2337 => x"ef004009",
        2338 => x"1305b400",
        2339 => x"93074400",
        2340 => x"137585ff",
        2341 => x"3307f540",
        2342 => x"e304f5f0",
        2343 => x"3304e400",
        2344 => x"b387a740",
        2345 => x"2320f400",
        2346 => x"6ff09fef",
        2347 => x"23a2e700",
        2348 => x"6ff05ffc",
        2349 => x"03274400",
        2350 => x"63968700",
        2351 => x"23a0e188",
        2352 => x"6ff01ffc",
        2353 => x"23a2e700",
        2354 => x"6ff09ffb",
        2355 => x"93070400",
        2356 => x"03244400",
        2357 => x"6ff0dfef",
        2358 => x"13840700",
        2359 => x"83a74700",
        2360 => x"6ff05ff1",
        2361 => x"13870700",
        2362 => x"83a74700",
        2363 => x"e39c87fe",
        2364 => x"23220700",
        2365 => x"6ff0dff8",
        2366 => x"9307c000",
        2367 => x"2320f900",
        2368 => x"13050900",
        2369 => x"ef004001",
        2370 => x"6ff05fe9",
        2371 => x"23209500",
        2372 => x"6ff01ff7",
        2373 => x"67800000",
        2374 => x"67800000",
        2375 => x"130101fe",
        2376 => x"23282101",
        2377 => x"03a98500",
        2378 => x"232c8100",
        2379 => x"23263101",
        2380 => x"23206101",
        2381 => x"232e1100",
        2382 => x"232a9100",
        2383 => x"23244101",
        2384 => x"23225101",
        2385 => x"13840500",
        2386 => x"130b0600",
        2387 => x"93890600",
        2388 => x"63ec2613",
        2389 => x"8397c500",
        2390 => x"13070900",
        2391 => x"93f60748",
        2392 => x"638c0608",
        2393 => x"83244401",
        2394 => x"13073000",
        2395 => x"83a50501",
        2396 => x"b384e402",
        2397 => x"13072000",
        2398 => x"032a0400",
        2399 => x"930a0500",
        2400 => x"330aba40",
        2401 => x"b3c4e402",
        2402 => x"13871900",
        2403 => x"33074701",
        2404 => x"13860400",
        2405 => x"63f6e400",
        2406 => x"93040700",
        2407 => x"13060700",
        2408 => x"93f70740",
        2409 => x"6386070a",
        2410 => x"93050600",
        2411 => x"13850a00",
        2412 => x"eff09fda",
        2413 => x"13090500",
        2414 => x"630a050a",
        2415 => x"83250401",
        2416 => x"13060a00",
        2417 => x"efe05fe1",
        2418 => x"8357c400",
        2419 => x"93f7f7b7",
        2420 => x"93e70708",
        2421 => x"2316f400",
        2422 => x"23282401",
        2423 => x"232a9400",
        2424 => x"33094901",
        2425 => x"b3844441",
        2426 => x"23202401",
        2427 => x"23249400",
        2428 => x"13890900",
        2429 => x"13870900",
        2430 => x"93090700",
        2431 => x"03250400",
        2432 => x"13860900",
        2433 => x"93050b00",
        2434 => x"efe05fdf",
        2435 => x"83278400",
        2436 => x"13050000",
        2437 => x"b3872741",
        2438 => x"2324f400",
        2439 => x"83270400",
        2440 => x"b3873701",
        2441 => x"2320f400",
        2442 => x"8320c101",
        2443 => x"03248101",
        2444 => x"83244101",
        2445 => x"03290101",
        2446 => x"8329c100",
        2447 => x"032a8100",
        2448 => x"832a4100",
        2449 => x"032b0100",
        2450 => x"13010102",
        2451 => x"67800000",
        2452 => x"13850a00",
        2453 => x"ef00105d",
        2454 => x"13090500",
        2455 => x"e31e05f6",
        2456 => x"83250401",
        2457 => x"13850a00",
        2458 => x"eff05fb7",
        2459 => x"9307c000",
        2460 => x"23a0fa00",
        2461 => x"8357c400",
        2462 => x"1305f0ff",
        2463 => x"93e70704",
        2464 => x"2316f400",
        2465 => x"6ff05ffa",
        2466 => x"13890600",
        2467 => x"6ff01ff7",
        2468 => x"83278600",
        2469 => x"130101fd",
        2470 => x"232e3101",
        2471 => x"23261102",
        2472 => x"23248102",
        2473 => x"23229102",
        2474 => x"23202103",
        2475 => x"232c4101",
        2476 => x"232a5101",
        2477 => x"23286101",
        2478 => x"23267101",
        2479 => x"23248101",
        2480 => x"23229101",
        2481 => x"2320a101",
        2482 => x"93090600",
        2483 => x"63800710",
        2484 => x"032a0600",
        2485 => x"930c0500",
        2486 => x"13840500",
        2487 => x"930a3000",
        2488 => x"130b2000",
        2489 => x"83270a00",
        2490 => x"032c4a00",
        2491 => x"138d0700",
        2492 => x"630e0c10",
        2493 => x"03298400",
        2494 => x"93040900",
        2495 => x"636a2c15",
        2496 => x"8317c400",
        2497 => x"13f70748",
        2498 => x"63060708",
        2499 => x"83244401",
        2500 => x"83250401",
        2501 => x"832b0400",
        2502 => x"b3845403",
        2503 => x"b38bbb40",
        2504 => x"13871b00",
        2505 => x"33078701",
        2506 => x"b3c46403",
        2507 => x"13860400",
        2508 => x"63f6e400",
        2509 => x"93040700",
        2510 => x"13060700",
        2511 => x"93f70740",
        2512 => x"638a070c",
        2513 => x"93050600",
        2514 => x"13850c00",
        2515 => x"eff0dfc0",
        2516 => x"13090500",
        2517 => x"630e050c",
        2518 => x"83250401",
        2519 => x"13860b00",
        2520 => x"efe09fc7",
        2521 => x"8357c400",
        2522 => x"93f7f7b7",
        2523 => x"93e70708",
        2524 => x"2316f400",
        2525 => x"23282401",
        2526 => x"232a9400",
        2527 => x"33097901",
        2528 => x"b3847441",
        2529 => x"23202401",
        2530 => x"23249400",
        2531 => x"13090c00",
        2532 => x"93040c00",
        2533 => x"03250400",
        2534 => x"13860400",
        2535 => x"93050d00",
        2536 => x"efe0dfc5",
        2537 => x"83278400",
        2538 => x"b3872741",
        2539 => x"2324f400",
        2540 => x"83270400",
        2541 => x"b3879700",
        2542 => x"2320f400",
        2543 => x"83a78900",
        2544 => x"b3878741",
        2545 => x"23a4f900",
        2546 => x"63920704",
        2547 => x"13050000",
        2548 => x"8320c102",
        2549 => x"03248102",
        2550 => x"23a20900",
        2551 => x"83244102",
        2552 => x"03290102",
        2553 => x"8329c101",
        2554 => x"032a8101",
        2555 => x"832a4101",
        2556 => x"032b0101",
        2557 => x"832bc100",
        2558 => x"032c8100",
        2559 => x"832c4100",
        2560 => x"032d0100",
        2561 => x"13010103",
        2562 => x"67800000",
        2563 => x"130a8a00",
        2564 => x"6ff05fed",
        2565 => x"13850c00",
        2566 => x"ef00d040",
        2567 => x"13090500",
        2568 => x"e31a05f4",
        2569 => x"83250401",
        2570 => x"13850c00",
        2571 => x"eff01f9b",
        2572 => x"9307c000",
        2573 => x"23a0fc00",
        2574 => x"8357c400",
        2575 => x"1305f0ff",
        2576 => x"93e70704",
        2577 => x"2316f400",
        2578 => x"23a40900",
        2579 => x"6ff05ff8",
        2580 => x"13090c00",
        2581 => x"6ff0dff3",
        2582 => x"83d7c500",
        2583 => x"130101f5",
        2584 => x"2322910a",
        2585 => x"23248109",
        2586 => x"2326110a",
        2587 => x"2324810a",
        2588 => x"2320210b",
        2589 => x"232e3109",
        2590 => x"232c4109",
        2591 => x"232a5109",
        2592 => x"23286109",
        2593 => x"23267109",
        2594 => x"93f70708",
        2595 => x"130c0500",
        2596 => x"93840500",
        2597 => x"638a0706",
        2598 => x"83a70501",
        2599 => x"63960706",
        2600 => x"93050004",
        2601 => x"2326d100",
        2602 => x"2324c100",
        2603 => x"eff0dfaa",
        2604 => x"23a0a400",
        2605 => x"23a8a400",
        2606 => x"03268100",
        2607 => x"8326c100",
        2608 => x"63100504",
        2609 => x"9307c000",
        2610 => x"2320fc00",
        2611 => x"1305f0ff",
        2612 => x"8320c10a",
        2613 => x"0324810a",
        2614 => x"8324410a",
        2615 => x"0329010a",
        2616 => x"8329c109",
        2617 => x"032a8109",
        2618 => x"832a4109",
        2619 => x"032b0109",
        2620 => x"832bc108",
        2621 => x"032c8108",
        2622 => x"1301010b",
        2623 => x"67800000",
        2624 => x"93070004",
        2625 => x"23aaf400",
        2626 => x"93070002",
        2627 => x"a30cf102",
        2628 => x"b7490000",
        2629 => x"93070003",
        2630 => x"232a0102",
        2631 => x"230df102",
        2632 => x"232ed100",
        2633 => x"130af0ff",
        2634 => x"938949b2",
        2635 => x"130b1000",
        2636 => x"930aa000",
        2637 => x"13040600",
        2638 => x"83470400",
        2639 => x"b33bf000",
        2640 => x"9387b7fd",
        2641 => x"b337f000",
        2642 => x"b3fbfb00",
        2643 => x"63900b0c",
        2644 => x"b306c440",
        2645 => x"6304c402",
        2646 => x"93850400",
        2647 => x"13050c00",
        2648 => x"2324d100",
        2649 => x"eff09fbb",
        2650 => x"630c4523",
        2651 => x"83274103",
        2652 => x"83268100",
        2653 => x"b387d700",
        2654 => x"232af102",
        2655 => x"83470400",
        2656 => x"63800722",
        2657 => x"13041400",
        2658 => x"23200102",
        2659 => x"23260102",
        2660 => x"23224103",
        2661 => x"23240102",
        2662 => x"a3010106",
        2663 => x"232c0106",
        2664 => x"83450400",
        2665 => x"13065000",
        2666 => x"13850900",
        2667 => x"ef00101c",
        2668 => x"83270102",
        2669 => x"93061400",
        2670 => x"631e0504",
        2671 => x"13f70701",
        2672 => x"63060700",
        2673 => x"13070002",
        2674 => x"a301e106",
        2675 => x"13f78700",
        2676 => x"63060700",
        2677 => x"1307b002",
        2678 => x"a301e106",
        2679 => x"03460400",
        2680 => x"1307a002",
        2681 => x"6304e604",
        2682 => x"8327c102",
        2683 => x"93060000",
        2684 => x"13069000",
        2685 => x"03470400",
        2686 => x"130707fd",
        2687 => x"637ee608",
        2688 => x"63840604",
        2689 => x"2326f102",
        2690 => x"6f000004",
        2691 => x"13041400",
        2692 => x"6ff09ff2",
        2693 => x"33053541",
        2694 => x"3315ab00",
        2695 => x"3365f500",
        2696 => x"2320a102",
        2697 => x"13840600",
        2698 => x"6ff09ff7",
        2699 => x"0327c101",
        2700 => x"13064700",
        2701 => x"03270700",
        2702 => x"232ec100",
        2703 => x"63440704",
        2704 => x"2326e102",
        2705 => x"13840600",
        2706 => x"03470400",
        2707 => x"9307e002",
        2708 => x"631ef706",
        2709 => x"03471400",
        2710 => x"9307a002",
        2711 => x"6318f704",
        2712 => x"8327c101",
        2713 => x"13042400",
        2714 => x"13874700",
        2715 => x"83a70700",
        2716 => x"232ee100",
        2717 => x"63d40700",
        2718 => x"9307f0ff",
        2719 => x"2322f102",
        2720 => x"6f00c004",
        2721 => x"3307e040",
        2722 => x"93e72700",
        2723 => x"2326e102",
        2724 => x"2320f102",
        2725 => x"6ff01ffb",
        2726 => x"b3875703",
        2727 => x"13041400",
        2728 => x"93061000",
        2729 => x"b387e700",
        2730 => x"6ff0dff4",
        2731 => x"13041400",
        2732 => x"23220102",
        2733 => x"93070000",
        2734 => x"93069000",
        2735 => x"03470400",
        2736 => x"130707fd",
        2737 => x"63f8e608",
        2738 => x"e39a0bfa",
        2739 => x"83450400",
        2740 => x"b74b0000",
        2741 => x"13063000",
        2742 => x"1385cbb2",
        2743 => x"ef001009",
        2744 => x"63020502",
        2745 => x"83270102",
        2746 => x"938bcbb2",
        2747 => x"33057541",
        2748 => x"13070004",
        2749 => x"3317a700",
        2750 => x"b3e7e700",
        2751 => x"13041400",
        2752 => x"2320f102",
        2753 => x"83450400",
        2754 => x"37450000",
        2755 => x"13066000",
        2756 => x"130505b3",
        2757 => x"230cb102",
        2758 => x"ef005005",
        2759 => x"630c0508",
        2760 => x"93070000",
        2761 => x"639a0704",
        2762 => x"03270102",
        2763 => x"8327c101",
        2764 => x"13770710",
        2765 => x"630a0702",
        2766 => x"93874700",
        2767 => x"232ef100",
        2768 => x"83274103",
        2769 => x"13061400",
        2770 => x"b3872701",
        2771 => x"232af102",
        2772 => x"6ff05fde",
        2773 => x"b3875703",
        2774 => x"13041400",
        2775 => x"930b1000",
        2776 => x"b387e700",
        2777 => x"6ff09ff5",
        2778 => x"93877700",
        2779 => x"93f787ff",
        2780 => x"93878700",
        2781 => x"6ff09ffc",
        2782 => x"b7260000",
        2783 => x"1307c101",
        2784 => x"9386c651",
        2785 => x"13860400",
        2786 => x"93050102",
        2787 => x"13050c00",
        2788 => x"97000000",
        2789 => x"e7000000",
        2790 => x"13090500",
        2791 => x"e31245fb",
        2792 => x"83d7c400",
        2793 => x"93f70704",
        2794 => x"e39207d2",
        2795 => x"03254103",
        2796 => x"6ff01fd2",
        2797 => x"b7260000",
        2798 => x"1307c101",
        2799 => x"9386c651",
        2800 => x"13860400",
        2801 => x"93050102",
        2802 => x"13050c00",
        2803 => x"ef00c01b",
        2804 => x"6ff09ffc",
        2805 => x"130101fd",
        2806 => x"232e3101",
        2807 => x"83a70501",
        2808 => x"93090700",
        2809 => x"03a78500",
        2810 => x"23248102",
        2811 => x"23202103",
        2812 => x"23286101",
        2813 => x"23267101",
        2814 => x"23261102",
        2815 => x"23229102",
        2816 => x"232c4101",
        2817 => x"232a5101",
        2818 => x"130b0500",
        2819 => x"13840500",
        2820 => x"13090600",
        2821 => x"938b0600",
        2822 => x"63d4e700",
        2823 => x"93070700",
        2824 => x"2320f900",
        2825 => x"03473404",
        2826 => x"63060700",
        2827 => x"93871700",
        2828 => x"2320f900",
        2829 => x"83270400",
        2830 => x"93f70702",
        2831 => x"63880700",
        2832 => x"83270900",
        2833 => x"93872700",
        2834 => x"2320f900",
        2835 => x"83240400",
        2836 => x"93f46400",
        2837 => x"639e0400",
        2838 => x"130a9401",
        2839 => x"930af0ff",
        2840 => x"8327c400",
        2841 => x"03270900",
        2842 => x"b387e740",
        2843 => x"63c4f408",
        2844 => x"83270400",
        2845 => x"83463404",
        2846 => x"93f70702",
        2847 => x"b336d000",
        2848 => x"6392070c",
        2849 => x"13063404",
        2850 => x"93850b00",
        2851 => x"13050b00",
        2852 => x"e7800900",
        2853 => x"9307f0ff",
        2854 => x"630af506",
        2855 => x"83270400",
        2856 => x"13074000",
        2857 => x"93040000",
        2858 => x"93f76700",
        2859 => x"639ee700",
        2860 => x"83270900",
        2861 => x"8324c400",
        2862 => x"b384f440",
        2863 => x"93c7f4ff",
        2864 => x"93d7f741",
        2865 => x"b3f4f400",
        2866 => x"83278400",
        2867 => x"03270401",
        2868 => x"6356f700",
        2869 => x"b387e740",
        2870 => x"b384f400",
        2871 => x"13090000",
        2872 => x"1304a401",
        2873 => x"130af0ff",
        2874 => x"63902409",
        2875 => x"13050000",
        2876 => x"6f000002",
        2877 => x"93061000",
        2878 => x"13060a00",
        2879 => x"93850b00",
        2880 => x"13050b00",
        2881 => x"e7800900",
        2882 => x"631a5503",
        2883 => x"1305f0ff",
        2884 => x"8320c102",
        2885 => x"03248102",
        2886 => x"83244102",
        2887 => x"03290102",
        2888 => x"8329c101",
        2889 => x"032a8101",
        2890 => x"832a4101",
        2891 => x"032b0101",
        2892 => x"832bc100",
        2893 => x"13010103",
        2894 => x"67800000",
        2895 => x"93841400",
        2896 => x"6ff01ff2",
        2897 => x"3307d400",
        2898 => x"13060003",
        2899 => x"a301c704",
        2900 => x"03475404",
        2901 => x"93871600",
        2902 => x"b307f400",
        2903 => x"93862600",
        2904 => x"a381e704",
        2905 => x"6ff01ff2",
        2906 => x"93061000",
        2907 => x"13060400",
        2908 => x"93850b00",
        2909 => x"13050b00",
        2910 => x"e7800900",
        2911 => x"e30845f9",
        2912 => x"13091900",
        2913 => x"6ff05ff6",
        2914 => x"130101fc",
        2915 => x"232c8102",
        2916 => x"232a9102",
        2917 => x"23244103",
        2918 => x"23225103",
        2919 => x"232e1102",
        2920 => x"23282103",
        2921 => x"23263103",
        2922 => x"83c78501",
        2923 => x"93840600",
        2924 => x"93068007",
        2925 => x"130a0500",
        2926 => x"13840500",
        2927 => x"930a0600",
        2928 => x"63eef600",
        2929 => x"93062006",
        2930 => x"13863504",
        2931 => x"63ecf600",
        2932 => x"63820728",
        2933 => x"93068005",
        2934 => x"638ed720",
        2935 => x"13092404",
        2936 => x"6f000004",
        2937 => x"9386d7f9",
        2938 => x"93f6f60f",
        2939 => x"93055001",
        2940 => x"e3e6d5fe",
        2941 => x"b7450000",
        2942 => x"93962600",
        2943 => x"938505b6",
        2944 => x"b386b600",
        2945 => x"83a60600",
        2946 => x"67800600",
        2947 => x"83270700",
        2948 => x"13092404",
        2949 => x"93864700",
        2950 => x"83a70700",
        2951 => x"2320d700",
        2952 => x"2301f404",
        2953 => x"93071000",
        2954 => x"6f008026",
        2955 => x"83270400",
        2956 => x"03250700",
        2957 => x"93f60708",
        2958 => x"93054500",
        2959 => x"63860602",
        2960 => x"83270500",
        2961 => x"2320b700",
        2962 => x"b7460000",
        2963 => x"63d80700",
        2964 => x"1307d002",
        2965 => x"b307f040",
        2966 => x"a301e404",
        2967 => x"938686b3",
        2968 => x"1307a000",
        2969 => x"6f008006",
        2970 => x"93f60704",
        2971 => x"83270500",
        2972 => x"2320b700",
        2973 => x"e38a06fc",
        2974 => x"93970701",
        2975 => x"93d70741",
        2976 => x"6ff09ffc",
        2977 => x"83250400",
        2978 => x"83260700",
        2979 => x"13f50508",
        2980 => x"83a70600",
        2981 => x"93864600",
        2982 => x"631a0500",
        2983 => x"93f50504",
        2984 => x"63860500",
        2985 => x"93970701",
        2986 => x"93d70701",
        2987 => x"2320d700",
        2988 => x"83458401",
        2989 => x"b7460000",
        2990 => x"1307f006",
        2991 => x"938686b3",
        2992 => x"6398e514",
        2993 => x"13078000",
        2994 => x"a3010404",
        2995 => x"83254400",
        2996 => x"2324b400",
        2997 => x"63ce0500",
        2998 => x"03250400",
        2999 => x"b3e5b700",
        3000 => x"13090600",
        3001 => x"1375b5ff",
        3002 => x"2320a400",
        3003 => x"63840502",
        3004 => x"13090600",
        3005 => x"b3f5e702",
        3006 => x"1309f9ff",
        3007 => x"b385b600",
        3008 => x"83c50500",
        3009 => x"2300b900",
        3010 => x"93850700",
        3011 => x"b3d7e702",
        3012 => x"e3f2e5fe",
        3013 => x"93078000",
        3014 => x"6314f702",
        3015 => x"83270400",
        3016 => x"93f71700",
        3017 => x"638e0700",
        3018 => x"03274400",
        3019 => x"83270401",
        3020 => x"63c8e700",
        3021 => x"93070003",
        3022 => x"a30ff9fe",
        3023 => x"1309f9ff",
        3024 => x"33062641",
        3025 => x"2328c400",
        3026 => x"13870400",
        3027 => x"93860a00",
        3028 => x"1306c101",
        3029 => x"93050400",
        3030 => x"13050a00",
        3031 => x"eff09fc7",
        3032 => x"9309f0ff",
        3033 => x"631c3513",
        3034 => x"1305f0ff",
        3035 => x"8320c103",
        3036 => x"03248103",
        3037 => x"83244103",
        3038 => x"03290103",
        3039 => x"8329c102",
        3040 => x"032a8102",
        3041 => x"832a4102",
        3042 => x"13010104",
        3043 => x"67800000",
        3044 => x"83270400",
        3045 => x"93e70702",
        3046 => x"2320f400",
        3047 => x"b7460000",
        3048 => x"93078007",
        3049 => x"9386c6b4",
        3050 => x"a302f404",
        3051 => x"83250400",
        3052 => x"03250700",
        3053 => x"13f80508",
        3054 => x"83270500",
        3055 => x"13054500",
        3056 => x"631a0800",
        3057 => x"13f80504",
        3058 => x"63060800",
        3059 => x"93970701",
        3060 => x"93d70701",
        3061 => x"2320a700",
        3062 => x"13f71500",
        3063 => x"63060700",
        3064 => x"93e50502",
        3065 => x"2320b400",
        3066 => x"638c0700",
        3067 => x"13070001",
        3068 => x"6ff09fed",
        3069 => x"b7460000",
        3070 => x"938686b3",
        3071 => x"6ff0dffa",
        3072 => x"03270400",
        3073 => x"1377f7fd",
        3074 => x"2320e400",
        3075 => x"6ff01ffe",
        3076 => x"1307a000",
        3077 => x"6ff05feb",
        3078 => x"83260400",
        3079 => x"83270700",
        3080 => x"83254401",
        3081 => x"13f80608",
        3082 => x"13854700",
        3083 => x"630a0800",
        3084 => x"2320a700",
        3085 => x"83a70700",
        3086 => x"23a0b700",
        3087 => x"6f008001",
        3088 => x"2320a700",
        3089 => x"93f60604",
        3090 => x"83a70700",
        3091 => x"e38606fe",
        3092 => x"2390b700",
        3093 => x"23280400",
        3094 => x"13090600",
        3095 => x"6ff0dfee",
        3096 => x"83270700",
        3097 => x"03264400",
        3098 => x"93050000",
        3099 => x"93864700",
        3100 => x"2320d700",
        3101 => x"03a90700",
        3102 => x"13050900",
        3103 => x"ef00002f",
        3104 => x"63060500",
        3105 => x"33052541",
        3106 => x"2322a400",
        3107 => x"83274400",
        3108 => x"2328f400",
        3109 => x"a3010404",
        3110 => x"6ff01feb",
        3111 => x"83260401",
        3112 => x"13060900",
        3113 => x"93850a00",
        3114 => x"13050a00",
        3115 => x"e7800400",
        3116 => x"e30c35eb",
        3117 => x"83270400",
        3118 => x"93f72700",
        3119 => x"63960704",
        3120 => x"8327c101",
        3121 => x"0325c400",
        3122 => x"e352f5ea",
        3123 => x"13850700",
        3124 => x"6ff0dfe9",
        3125 => x"93061000",
        3126 => x"93850a00",
        3127 => x"13050a00",
        3128 => x"2326c100",
        3129 => x"e7800400",
        3130 => x"e30035e9",
        3131 => x"0326c100",
        3132 => x"13091900",
        3133 => x"8327c400",
        3134 => x"0327c101",
        3135 => x"b387e740",
        3136 => x"e34af9fc",
        3137 => x"6ff0dffb",
        3138 => x"13090000",
        3139 => x"13069401",
        3140 => x"6ff05ffe",
        3141 => x"8397c500",
        3142 => x"130101fe",
        3143 => x"232c8100",
        3144 => x"232a9100",
        3145 => x"232e1100",
        3146 => x"23282101",
        3147 => x"13f78700",
        3148 => x"93040500",
        3149 => x"13840500",
        3150 => x"63120712",
        3151 => x"03a74500",
        3152 => x"6346e000",
        3153 => x"03a70504",
        3154 => x"6356e010",
        3155 => x"0327c402",
        3156 => x"63020710",
        3157 => x"03a90400",
        3158 => x"93963701",
        3159 => x"23a00400",
        3160 => x"63dc060a",
        3161 => x"03264405",
        3162 => x"8357c400",
        3163 => x"93f74700",
        3164 => x"638e0700",
        3165 => x"83274400",
        3166 => x"3306f640",
        3167 => x"83274403",
        3168 => x"63860700",
        3169 => x"83270404",
        3170 => x"3306f640",
        3171 => x"8327c402",
        3172 => x"83250402",
        3173 => x"93060000",
        3174 => x"13850400",
        3175 => x"e7800700",
        3176 => x"1307f0ff",
        3177 => x"8317c400",
        3178 => x"6312e502",
        3179 => x"83a60400",
        3180 => x"1307d001",
        3181 => x"636cd70e",
        3182 => x"37074020",
        3183 => x"13071700",
        3184 => x"3357d700",
        3185 => x"13771700",
        3186 => x"6302070e",
        3187 => x"03270401",
        3188 => x"23220400",
        3189 => x"2320e400",
        3190 => x"13973701",
        3191 => x"635c0700",
        3192 => x"9307f0ff",
        3193 => x"6316f500",
        3194 => x"83a70400",
        3195 => x"63940700",
        3196 => x"232aa404",
        3197 => x"83254403",
        3198 => x"23a02401",
        3199 => x"638c0504",
        3200 => x"93074404",
        3201 => x"6386f500",
        3202 => x"13850400",
        3203 => x"efe01ffd",
        3204 => x"232a0402",
        3205 => x"6f000004",
        3206 => x"83250402",
        3207 => x"13060000",
        3208 => x"93061000",
        3209 => x"13850400",
        3210 => x"e7000700",
        3211 => x"9307f0ff",
        3212 => x"13060500",
        3213 => x"e31af5f2",
        3214 => x"83a70400",
        3215 => x"e38607f2",
        3216 => x"138737fe",
        3217 => x"63060700",
        3218 => x"9387a7fe",
        3219 => x"639e0704",
        3220 => x"23a02401",
        3221 => x"13050000",
        3222 => x"6f000006",
        3223 => x"03a60501",
        3224 => x"e30a06fe",
        3225 => x"83a60500",
        3226 => x"93f73700",
        3227 => x"23a0c500",
        3228 => x"3389c640",
        3229 => x"13070000",
        3230 => x"63940700",
        3231 => x"03a74501",
        3232 => x"2324e400",
        3233 => x"e35820fd",
        3234 => x"83278402",
        3235 => x"83250402",
        3236 => x"93060900",
        3237 => x"13850400",
        3238 => x"2326c100",
        3239 => x"e7800700",
        3240 => x"0326c100",
        3241 => x"6346a002",
        3242 => x"8357c400",
        3243 => x"93e70704",
        3244 => x"2316f400",
        3245 => x"1305f0ff",
        3246 => x"8320c101",
        3247 => x"03248101",
        3248 => x"83244101",
        3249 => x"03290101",
        3250 => x"13010102",
        3251 => x"67800000",
        3252 => x"3306a600",
        3253 => x"3309a940",
        3254 => x"6ff0dffa",
        3255 => x"83a70501",
        3256 => x"638e0704",
        3257 => x"130101fe",
        3258 => x"232c8100",
        3259 => x"232e1100",
        3260 => x"13040500",
        3261 => x"630c0500",
        3262 => x"83270502",
        3263 => x"63980700",
        3264 => x"2326b100",
        3265 => x"efe09f86",
        3266 => x"8325c100",
        3267 => x"8397c500",
        3268 => x"638c0700",
        3269 => x"13050400",
        3270 => x"03248101",
        3271 => x"8320c101",
        3272 => x"13010102",
        3273 => x"6ff01fdf",
        3274 => x"8320c101",
        3275 => x"03248101",
        3276 => x"13050000",
        3277 => x"13010102",
        3278 => x"67800000",
        3279 => x"13050000",
        3280 => x"67800000",
        3281 => x"93050500",
        3282 => x"631e0500",
        3283 => x"b7350000",
        3284 => x"37050020",
        3285 => x"13868181",
        3286 => x"9385c52d",
        3287 => x"13054502",
        3288 => x"6fe01f86",
        3289 => x"03a50187",
        3290 => x"6ff05ff7",
        3291 => x"93f5f50f",
        3292 => x"3306c500",
        3293 => x"6316c500",
        3294 => x"13050000",
        3295 => x"67800000",
        3296 => x"83470500",
        3297 => x"e38cb7fe",
        3298 => x"13051500",
        3299 => x"6ff09ffe",
        3300 => x"130101ff",
        3301 => x"23248100",
        3302 => x"23229100",
        3303 => x"93040500",
        3304 => x"13850500",
        3305 => x"93050600",
        3306 => x"23261100",
        3307 => x"23ac0186",
        3308 => x"ef00c01b",
        3309 => x"9307f0ff",
        3310 => x"6318f500",
        3311 => x"83a78187",
        3312 => x"63840700",
        3313 => x"23a0f400",
        3314 => x"8320c100",
        3315 => x"03248100",
        3316 => x"83244100",
        3317 => x"13010101",
        3318 => x"67800000",
        3319 => x"130101ff",
        3320 => x"23248100",
        3321 => x"23229100",
        3322 => x"93040500",
        3323 => x"13850500",
        3324 => x"23261100",
        3325 => x"23ac0186",
        3326 => x"ef008026",
        3327 => x"9307f0ff",
        3328 => x"6318f500",
        3329 => x"83a78187",
        3330 => x"63840700",
        3331 => x"23a0f400",
        3332 => x"8320c100",
        3333 => x"03248100",
        3334 => x"83244100",
        3335 => x"13010101",
        3336 => x"67800000",
        3337 => x"63960500",
        3338 => x"93050600",
        3339 => x"6fe0dff2",
        3340 => x"130101fe",
        3341 => x"232c8100",
        3342 => x"23244101",
        3343 => x"232e1100",
        3344 => x"232a9100",
        3345 => x"23282101",
        3346 => x"23263101",
        3347 => x"13040600",
        3348 => x"130a0500",
        3349 => x"63180602",
        3350 => x"efe05fd8",
        3351 => x"93040000",
        3352 => x"8320c101",
        3353 => x"03248101",
        3354 => x"03290101",
        3355 => x"8329c100",
        3356 => x"032a8100",
        3357 => x"13850400",
        3358 => x"83244101",
        3359 => x"13010102",
        3360 => x"67800000",
        3361 => x"93840500",
        3362 => x"ef008005",
        3363 => x"13090500",
        3364 => x"63668500",
        3365 => x"93571500",
        3366 => x"e3e487fc",
        3367 => x"93050400",
        3368 => x"13050a00",
        3369 => x"efe05feb",
        3370 => x"93090500",
        3371 => x"63160500",
        3372 => x"93840900",
        3373 => x"6ff0dffa",
        3374 => x"13060400",
        3375 => x"63748900",
        3376 => x"13060900",
        3377 => x"93850400",
        3378 => x"13850900",
        3379 => x"efd0dff0",
        3380 => x"93850400",
        3381 => x"13050a00",
        3382 => x"efe05fd0",
        3383 => x"6ff05ffd",
        3384 => x"83a7c5ff",
        3385 => x"1385c7ff",
        3386 => x"63d80700",
        3387 => x"b385a500",
        3388 => x"83a70500",
        3389 => x"3305f500",
        3390 => x"67800000",
        3391 => x"130101ff",
        3392 => x"23261100",
        3393 => x"23248100",
        3394 => x"93089003",
        3395 => x"73000000",
        3396 => x"13040500",
        3397 => x"635a0500",
        3398 => x"33048040",
        3399 => x"efe05fc1",
        3400 => x"23208500",
        3401 => x"1304f0ff",
        3402 => x"8320c100",
        3403 => x"13050400",
        3404 => x"03248100",
        3405 => x"13010101",
        3406 => x"67800000",
        3407 => x"9308d005",
        3408 => x"73000000",
        3409 => x"63520502",
        3410 => x"130101ff",
        3411 => x"23248100",
        3412 => x"13040500",
        3413 => x"23261100",
        3414 => x"33048040",
        3415 => x"efe05fbd",
        3416 => x"23208500",
        3417 => x"6f000000",
        3418 => x"6f000000",
        3419 => x"130101fe",
        3420 => x"232a9100",
        3421 => x"232e1100",
        3422 => x"93040500",
        3423 => x"232c8100",
        3424 => x"93083019",
        3425 => x"13050000",
        3426 => x"93050100",
        3427 => x"73000000",
        3428 => x"13040500",
        3429 => x"635a0500",
        3430 => x"33048040",
        3431 => x"efe05fb9",
        3432 => x"23208500",
        3433 => x"1304f0ff",
        3434 => x"83274100",
        3435 => x"03270100",
        3436 => x"8320c101",
        3437 => x"23a2f400",
        3438 => x"83278100",
        3439 => x"23a0e400",
        3440 => x"1307803e",
        3441 => x"b3c7e702",
        3442 => x"13050400",
        3443 => x"03248101",
        3444 => x"23a4f400",
        3445 => x"83244101",
        3446 => x"13010102",
        3447 => x"67800000",
        3448 => x"130101ff",
        3449 => x"23261100",
        3450 => x"23248100",
        3451 => x"9308e003",
        3452 => x"73000000",
        3453 => x"13040500",
        3454 => x"635a0500",
        3455 => x"33048040",
        3456 => x"efe01fb3",
        3457 => x"23208500",
        3458 => x"1304f0ff",
        3459 => x"8320c100",
        3460 => x"13050400",
        3461 => x"03248100",
        3462 => x"13010101",
        3463 => x"67800000",
        3464 => x"130101ff",
        3465 => x"23261100",
        3466 => x"23248100",
        3467 => x"9308f003",
        3468 => x"73000000",
        3469 => x"13040500",
        3470 => x"635a0500",
        3471 => x"33048040",
        3472 => x"efe01faf",
        3473 => x"23208500",
        3474 => x"1304f0ff",
        3475 => x"8320c100",
        3476 => x"13050400",
        3477 => x"03248100",
        3478 => x"13010101",
        3479 => x"67800000",
        3480 => x"93060500",
        3481 => x"03a54188",
        3482 => x"130101ff",
        3483 => x"23261100",
        3484 => x"631a0502",
        3485 => x"9308600d",
        3486 => x"73000000",
        3487 => x"9307f0ff",
        3488 => x"6310f502",
        3489 => x"efe0dfaa",
        3490 => x"9307c000",
        3491 => x"2320f500",
        3492 => x"1305f0ff",
        3493 => x"8320c100",
        3494 => x"13010101",
        3495 => x"67800000",
        3496 => x"23a2a188",
        3497 => x"9308600d",
        3498 => x"3385a600",
        3499 => x"73000000",
        3500 => x"83a74188",
        3501 => x"b386f600",
        3502 => x"e316d5fc",
        3503 => x"23a2a188",
        3504 => x"13850700",
        3505 => x"6ff01ffd",
        3506 => x"130101ff",
        3507 => x"23261100",
        3508 => x"23248100",
        3509 => x"93080004",
        3510 => x"73000000",
        3511 => x"13040500",
        3512 => x"635a0500",
        3513 => x"33048040",
        3514 => x"efe09fa4",
        3515 => x"23208500",
        3516 => x"1304f0ff",
        3517 => x"8320c100",
        3518 => x"13050400",
        3519 => x"03248100",
        3520 => x"13010101",
        3521 => x"67800000",
        3522 => x"10000000",
        3523 => x"00000000",
        3524 => x"037a5200",
        3525 => x"017c0101",
        3526 => x"1b0c0200",
        3527 => x"10000000",
        3528 => x"18000000",
        3529 => x"84d0ffff",
        3530 => x"0c040000",
        3531 => x"00000000",
        3532 => x"10000000",
        3533 => x"00000000",
        3534 => x"037a5200",
        3535 => x"017c0101",
        3536 => x"1b0c0200",
        3537 => x"10000000",
        3538 => x"18000000",
        3539 => x"68d4ffff",
        3540 => x"ec030000",
        3541 => x"00000000",
        3542 => x"10000000",
        3543 => x"00000000",
        3544 => x"037a5200",
        3545 => x"017c0101",
        3546 => x"1b0c0200",
        3547 => x"10000000",
        3548 => x"18000000",
        3549 => x"2cd8ffff",
        3550 => x"1c040000",
        3551 => x"00000000",
        3552 => x"30313233",
        3553 => x"34353637",
        3554 => x"38396162",
        3555 => x"63646566",
        3556 => x"00000000",
        3557 => x"a0040000",
        3558 => x"a4040000",
        3559 => x"a4040000",
        3560 => x"a4040000",
        3561 => x"14050000",
        3562 => x"a4040000",
        3563 => x"a4040000",
        3564 => x"a4040000",
        3565 => x"a4040000",
        3566 => x"a4040000",
        3567 => x"a4040000",
        3568 => x"a4040000",
        3569 => x"a4040000",
        3570 => x"a4040000",
        3571 => x"a4040000",
        3572 => x"1c050000",
        3573 => x"a4040000",
        3574 => x"34050000",
        3575 => x"3c050000",
        3576 => x"a4040000",
        3577 => x"44050000",
        3578 => x"4c050000",
        3579 => x"a4040000",
        3580 => x"24050000",
        3581 => x"2c050000",
        3582 => x"ac050000",
        3583 => x"80050000",
        3584 => x"80050000",
        3585 => x"80050000",
        3586 => x"80050000",
        3587 => x"a4040000",
        3588 => x"30060000",
        3589 => x"fc050000",
        3590 => x"80050000",
        3591 => x"80050000",
        3592 => x"80050000",
        3593 => x"80050000",
        3594 => x"80050000",
        3595 => x"80050000",
        3596 => x"80050000",
        3597 => x"80050000",
        3598 => x"80050000",
        3599 => x"80050000",
        3600 => x"80050000",
        3601 => x"80050000",
        3602 => x"80050000",
        3603 => x"80050000",
        3604 => x"a0050000",
        3605 => x"a0050000",
        3606 => x"80050000",
        3607 => x"80050000",
        3608 => x"80050000",
        3609 => x"80050000",
        3610 => x"80050000",
        3611 => x"80050000",
        3612 => x"80050000",
        3613 => x"80050000",
        3614 => x"80050000",
        3615 => x"80050000",
        3616 => x"80050000",
        3617 => x"80050000",
        3618 => x"a4040000",
        3619 => x"ac050000",
        3620 => x"c0050000",
        3621 => x"e8050000",
        3622 => x"80050000",
        3623 => x"80050000",
        3624 => x"80050000",
        3625 => x"80050000",
        3626 => x"80050000",
        3627 => x"80050000",
        3628 => x"d4050000",
        3629 => x"80050000",
        3630 => x"80050000",
        3631 => x"80050000",
        3632 => x"80050000",
        3633 => x"94050000",
        3634 => x"a0050000",
        3635 => x"00010202",
        3636 => x"03030303",
        3637 => x"04040404",
        3638 => x"04040404",
        3639 => x"05050505",
        3640 => x"05050505",
        3641 => x"05050505",
        3642 => x"05050505",
        3643 => x"06060606",
        3644 => x"06060606",
        3645 => x"06060606",
        3646 => x"06060606",
        3647 => x"06060606",
        3648 => x"06060606",
        3649 => x"06060606",
        3650 => x"06060606",
        3651 => x"07070707",
        3652 => x"07070707",
        3653 => x"07070707",
        3654 => x"07070707",
        3655 => x"07070707",
        3656 => x"07070707",
        3657 => x"07070707",
        3658 => x"07070707",
        3659 => x"07070707",
        3660 => x"07070707",
        3661 => x"07070707",
        3662 => x"07070707",
        3663 => x"07070707",
        3664 => x"07070707",
        3665 => x"07070707",
        3666 => x"07070707",
        3667 => x"08080808",
        3668 => x"08080808",
        3669 => x"08080808",
        3670 => x"08080808",
        3671 => x"08080808",
        3672 => x"08080808",
        3673 => x"08080808",
        3674 => x"08080808",
        3675 => x"08080808",
        3676 => x"08080808",
        3677 => x"08080808",
        3678 => x"08080808",
        3679 => x"08080808",
        3680 => x"08080808",
        3681 => x"08080808",
        3682 => x"08080808",
        3683 => x"08080808",
        3684 => x"08080808",
        3685 => x"08080808",
        3686 => x"08080808",
        3687 => x"08080808",
        3688 => x"08080808",
        3689 => x"08080808",
        3690 => x"08080808",
        3691 => x"08080808",
        3692 => x"08080808",
        3693 => x"08080808",
        3694 => x"08080808",
        3695 => x"08080808",
        3696 => x"08080808",
        3697 => x"08080808",
        3698 => x"08080808",
        3699 => x"0d0a4542",
        3700 => x"5245414b",
        3701 => x"21206d65",
        3702 => x"7063203d",
        3703 => x"20000000",
        3704 => x"20696e73",
        3705 => x"6e203d20",
        3706 => x"00000000",
        3707 => x"0d0a0000",
        3708 => x"0d0a0a44",
        3709 => x"6973706c",
        3710 => x"6179696e",
        3711 => x"67207468",
        3712 => x"65207469",
        3713 => x"6d652070",
        3714 => x"61737365",
        3715 => x"64207369",
        3716 => x"6e636520",
        3717 => x"72657365",
        3718 => x"740d0a0a",
        3719 => x"00000000",
        3720 => x"4f6e2d63",
        3721 => x"68697020",
        3722 => x"64656275",
        3723 => x"67676572",
        3724 => x"20666f75",
        3725 => x"6e642c20",
        3726 => x"736b6970",
        3727 => x"70696e67",
        3728 => x"20454252",
        3729 => x"45414b20",
        3730 => x"696e7374",
        3731 => x"72756374",
        3732 => x"696f6e0d",
        3733 => x"0a0d0a00",
        3734 => x"2530356c",
        3735 => x"643a2530",
        3736 => x"366c6420",
        3737 => x"20202530",
        3738 => x"326c643a",
        3739 => x"2530326c",
        3740 => x"643a2530",
        3741 => x"326c640d",
        3742 => x"00000000",
        3743 => x"696e7465",
        3744 => x"72727570",
        3745 => x"745f6469",
        3746 => x"72656374",
        3747 => x"00000000",
        3748 => x"54485541",
        3749 => x"53205249",
        3750 => x"53432d56",
        3751 => x"20525633",
        3752 => x"32494d20",
        3753 => x"62617265",
        3754 => x"206d6574",
        3755 => x"616c2070",
        3756 => x"726f6365",
        3757 => x"73736f72",
        3758 => x"00000000",
        3759 => x"54686520",
        3760 => x"48616775",
        3761 => x"6520556e",
        3762 => x"69766572",
        3763 => x"73697479",
        3764 => x"206f6620",
        3765 => x"4170706c",
        3766 => x"69656420",
        3767 => x"53636965",
        3768 => x"6e636573",
        3769 => x"00000000",
        3770 => x"44657061",
        3771 => x"72746d65",
        3772 => x"6e74206f",
        3773 => x"6620456c",
        3774 => x"65637472",
        3775 => x"6963616c",
        3776 => x"20456e67",
        3777 => x"696e6565",
        3778 => x"72696e67",
        3779 => x"00000000",
        3780 => x"4a2e452e",
        3781 => x"4a2e206f",
        3782 => x"70206465",
        3783 => x"6e204272",
        3784 => x"6f757700",
        3785 => x"232d302b",
        3786 => x"20000000",
        3787 => x"686c4c00",
        3788 => x"65666745",
        3789 => x"46470000",
        3790 => x"30313233",
        3791 => x"34353637",
        3792 => x"38394142",
        3793 => x"43444546",
        3794 => x"00000000",
        3795 => x"30313233",
        3796 => x"34353637",
        3797 => x"38396162",
        3798 => x"63646566",
        3799 => x"00000000",
        3800 => x"0c2e0000",
        3801 => x"2c2e0000",
        3802 => x"dc2d0000",
        3803 => x"dc2d0000",
        3804 => x"dc2d0000",
        3805 => x"dc2d0000",
        3806 => x"2c2e0000",
        3807 => x"dc2d0000",
        3808 => x"dc2d0000",
        3809 => x"dc2d0000",
        3810 => x"dc2d0000",
        3811 => x"18300000",
        3812 => x"842e0000",
        3813 => x"902f0000",
        3814 => x"dc2d0000",
        3815 => x"dc2d0000",
        3816 => x"60300000",
        3817 => x"dc2d0000",
        3818 => x"842e0000",
        3819 => x"dc2d0000",
        3820 => x"dc2d0000",
        3821 => x"9c2f0000",
        3822 => x"7c3a0000",
        3823 => x"903a0000",
        3824 => x"bc3a0000",
        3825 => x"e83a0000",
        3826 => x"103b0000",
        3827 => x"00000000",
        3828 => x"00000000",
        3829 => x"03000000",
        3830 => x"88000020",
        3831 => x"00000000",
        3832 => x"88000020",
        3833 => x"f0000020",
        3834 => x"58010020",
        3835 => x"00000000",
        3836 => x"00000000",
        3837 => x"00000000",
        3838 => x"00000000",
        3839 => x"00000000",
        3840 => x"00000000",
        3841 => x"00000000",
        3842 => x"00000000",
        3843 => x"00000000",
        3844 => x"00000000",
        3845 => x"00000000",
        3846 => x"00000000",
        3847 => x"00000000",
        3848 => x"00000000",
        3849 => x"00000000",
        3850 => x"24000020"
            );
end package rom_image;
