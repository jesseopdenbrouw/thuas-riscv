-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Sun Feb 25 19:27:05 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382022f",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"13868187",
           8 => x"9387819c",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13858187",
          13 => x"ef104035",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93878187",
          17 => x"637cf600",
          18 => x"b7450000",
          19 => x"3386c740",
          20 => x"938505c4",
          21 => x"13050500",
          22 => x"ef10c034",
          23 => x"ef208032",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef108072",
          29 => x"ef10102c",
          30 => x"6f104067",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef10406b",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"232c4101",
          40 => x"130a0500",
          41 => x"37450000",
          42 => x"1305c5a8",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"13044100",
          50 => x"ef100069",
          51 => x"37490000",
          52 => x"9309c1ff",
          53 => x"93070400",
          54 => x"13090981",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef108065",
          65 => x"37450000",
          66 => x"130505aa",
          67 => x"ef10c064",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef104062",
          78 => x"37450000",
          79 => x"1305c5aa",
          80 => x"ef108061",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74708",
          91 => x"b70600f0",
          92 => x"1377f7fe",
          93 => x"23a2e708",
          94 => x"83a74600",
          95 => x"93c71700",
          96 => x"23a2f600",
          97 => x"67800000",
          98 => x"370700f0",
          99 => x"83274700",
         100 => x"93e70720",
         101 => x"2322f700",
         102 => x"6f000000",
         103 => x"b70700f0",
         104 => x"b70500f0",
         105 => x"370500f0",
         106 => x"9387470f",
         107 => x"9385050f",
         108 => x"83a60700",
         109 => x"03a60500",
         110 => x"03a70700",
         111 => x"e31ad7fe",
         112 => x"b7870100",
         113 => x"b70500f0",
         114 => x"1308f0ff",
         115 => x"9387076a",
         116 => x"23ae050f",
         117 => x"b307f600",
         118 => x"b70600f0",
         119 => x"23ac060f",
         120 => x"33b6c700",
         121 => x"23acf60e",
         122 => x"3306e600",
         123 => x"23aec50e",
         124 => x"83274500",
         125 => x"93c72700",
         126 => x"2322f500",
         127 => x"67800000",
         128 => x"b70700f0",
         129 => x"03a74702",
         130 => x"b70600f0",
         131 => x"93870702",
         132 => x"13774700",
         133 => x"630a0700",
         134 => x"03a74600",
         135 => x"13478700",
         136 => x"23a2e600",
         137 => x"83a78700",
         138 => x"67800000",
         139 => x"b70700f0",
         140 => x"03a7470a",
         141 => x"b70600f0",
         142 => x"1377f7f0",
         143 => x"23a2e70a",
         144 => x"83a74600",
         145 => x"93c74700",
         146 => x"23a2f600",
         147 => x"67800000",
         148 => x"b70700f0",
         149 => x"03a74706",
         150 => x"b70600f0",
         151 => x"137777ff",
         152 => x"23a2e706",
         153 => x"83a74600",
         154 => x"93c70701",
         155 => x"23a2f600",
         156 => x"67800000",
         157 => x"b70700f0",
         158 => x"03a74704",
         159 => x"b70600f0",
         160 => x"137777ff",
         161 => x"23a2e704",
         162 => x"83a74600",
         163 => x"93c70702",
         164 => x"23a2f600",
         165 => x"67800000",
         166 => x"b70700f0",
         167 => x"03a74705",
         168 => x"b70600f0",
         169 => x"137777ff",
         170 => x"23aae704",
         171 => x"83a74600",
         172 => x"93c70708",
         173 => x"23a2f600",
         174 => x"67800000",
         175 => x"b70700f0",
         176 => x"23ae0700",
         177 => x"03a74700",
         178 => x"13470704",
         179 => x"23a2e700",
         180 => x"67800000",
         181 => x"370700f0",
         182 => x"b70600f0",
         183 => x"2326070e",
         184 => x"83a74600",
         185 => x"93c70710",
         186 => x"23a2f600",
         187 => x"67800000",
         188 => x"6f000000",
         189 => x"13050000",
         190 => x"67800000",
         191 => x"13050000",
         192 => x"67800000",
         193 => x"130101f7",
         194 => x"23221100",
         195 => x"23242100",
         196 => x"23263100",
         197 => x"23284100",
         198 => x"232a5100",
         199 => x"232c6100",
         200 => x"232e7100",
         201 => x"23208102",
         202 => x"23229102",
         203 => x"2324a102",
         204 => x"2326b102",
         205 => x"2328c102",
         206 => x"232ad102",
         207 => x"232ce102",
         208 => x"232ef102",
         209 => x"23200105",
         210 => x"23221105",
         211 => x"23242105",
         212 => x"23263105",
         213 => x"23284105",
         214 => x"232a5105",
         215 => x"232c6105",
         216 => x"232e7105",
         217 => x"23208107",
         218 => x"23229107",
         219 => x"2324a107",
         220 => x"2326b107",
         221 => x"2328c107",
         222 => x"232ad107",
         223 => x"232ce107",
         224 => x"232ef107",
         225 => x"f3222034",
         226 => x"23205108",
         227 => x"f3221034",
         228 => x"23225108",
         229 => x"83a20200",
         230 => x"23245108",
         231 => x"f3223034",
         232 => x"23265108",
         233 => x"f3272034",
         234 => x"1307b000",
         235 => x"6374f70c",
         236 => x"37070080",
         237 => x"1307d7ff",
         238 => x"b387e700",
         239 => x"13078001",
         240 => x"636ef700",
         241 => x"37470000",
         242 => x"93972700",
         243 => x"13074782",
         244 => x"b387e700",
         245 => x"83a70700",
         246 => x"67800700",
         247 => x"03258102",
         248 => x"83220108",
         249 => x"63c80200",
         250 => x"f3221034",
         251 => x"93824200",
         252 => x"73901234",
         253 => x"832fc107",
         254 => x"032f8107",
         255 => x"832e4107",
         256 => x"032e0107",
         257 => x"832dc106",
         258 => x"032d8106",
         259 => x"832c4106",
         260 => x"032c0106",
         261 => x"832bc105",
         262 => x"032b8105",
         263 => x"832a4105",
         264 => x"032a0105",
         265 => x"8329c104",
         266 => x"03298104",
         267 => x"83284104",
         268 => x"03280104",
         269 => x"8327c103",
         270 => x"03278103",
         271 => x"83264103",
         272 => x"03260103",
         273 => x"8325c102",
         274 => x"83244102",
         275 => x"03240102",
         276 => x"8323c101",
         277 => x"03238101",
         278 => x"83224101",
         279 => x"03220101",
         280 => x"8321c100",
         281 => x"03218100",
         282 => x"83204100",
         283 => x"13010109",
         284 => x"73002030",
         285 => x"93061000",
         286 => x"e3f2f6f6",
         287 => x"e360f7f6",
         288 => x"37470000",
         289 => x"93972700",
         290 => x"13078788",
         291 => x"b387e700",
         292 => x"83a70700",
         293 => x"67800700",
         294 => x"eff09fdb",
         295 => x"03258102",
         296 => x"6ff01ff4",
         297 => x"eff01fe3",
         298 => x"03258102",
         299 => x"6ff05ff3",
         300 => x"eff0dfce",
         301 => x"03258102",
         302 => x"6ff09ff2",
         303 => x"eff01fe0",
         304 => x"03258102",
         305 => x"6ff0dff1",
         306 => x"eff0dfc9",
         307 => x"03258102",
         308 => x"6ff01ff1",
         309 => x"eff09fd5",
         310 => x"03258102",
         311 => x"6ff05ff0",
         312 => x"eff01fd2",
         313 => x"03258102",
         314 => x"6ff09fef",
         315 => x"eff0dfda",
         316 => x"03258102",
         317 => x"6ff0dfee",
         318 => x"eff0dfd7",
         319 => x"03258102",
         320 => x"6ff01fee",
         321 => x"13050100",
         322 => x"eff01fb9",
         323 => x"03258102",
         324 => x"6ff01fed",
         325 => x"9307900a",
         326 => x"6380f814",
         327 => x"63d81703",
         328 => x"9307600d",
         329 => x"638ef818",
         330 => x"938808c0",
         331 => x"9307f000",
         332 => x"63e01705",
         333 => x"b7470000",
         334 => x"9387878b",
         335 => x"93982800",
         336 => x"b388f800",
         337 => x"83a70800",
         338 => x"67800700",
         339 => x"938878fc",
         340 => x"93074002",
         341 => x"63ee1701",
         342 => x"b7470000",
         343 => x"9387878f",
         344 => x"93982800",
         345 => x"b388f800",
         346 => x"83a70800",
         347 => x"67800700",
         348 => x"ef10d060",
         349 => x"93078005",
         350 => x"2320f500",
         351 => x"9307f0ff",
         352 => x"13850700",
         353 => x"6ff0dfe5",
         354 => x"b7270000",
         355 => x"23a2f500",
         356 => x"93070000",
         357 => x"13850700",
         358 => x"6ff09fe4",
         359 => x"93070000",
         360 => x"13850700",
         361 => x"6ff0dfe3",
         362 => x"ef10505d",
         363 => x"93079000",
         364 => x"2320f500",
         365 => x"9307f0ff",
         366 => x"13850700",
         367 => x"6ff05fe2",
         368 => x"ef10d05b",
         369 => x"9307f001",
         370 => x"2320f500",
         371 => x"9307f0ff",
         372 => x"13850700",
         373 => x"6ff0dfe0",
         374 => x"ef10505a",
         375 => x"9307d000",
         376 => x"2320f500",
         377 => x"9307f0ff",
         378 => x"13850700",
         379 => x"6ff05fdf",
         380 => x"ef10d058",
         381 => x"93072000",
         382 => x"2320f500",
         383 => x"9307f0ff",
         384 => x"13850700",
         385 => x"6ff0dfdd",
         386 => x"13090600",
         387 => x"13840500",
         388 => x"635cc000",
         389 => x"b384c500",
         390 => x"eff01fa6",
         391 => x"2300a400",
         392 => x"13041400",
         393 => x"e39a84fe",
         394 => x"13050900",
         395 => x"6ff05fdb",
         396 => x"13090600",
         397 => x"13840500",
         398 => x"e358c0fe",
         399 => x"b384c500",
         400 => x"03450400",
         401 => x"13041400",
         402 => x"eff05fa3",
         403 => x"e39a84fe",
         404 => x"13050900",
         405 => x"6ff0dfd8",
         406 => x"13090000",
         407 => x"93040500",
         408 => x"13040900",
         409 => x"93090900",
         410 => x"93070900",
         411 => x"732410c8",
         412 => x"f32910c0",
         413 => x"f32710c8",
         414 => x"e31af4fe",
         415 => x"37460f00",
         416 => x"13060624",
         417 => x"93060000",
         418 => x"13850900",
         419 => x"93050400",
         420 => x"ef005011",
         421 => x"37460f00",
         422 => x"23a4a400",
         423 => x"13060624",
         424 => x"93060000",
         425 => x"13850900",
         426 => x"93050400",
         427 => x"ef00804c",
         428 => x"23a0a400",
         429 => x"23a2b400",
         430 => x"13050900",
         431 => x"6ff05fd2",
         432 => x"63180500",
         433 => x"1385819c",
         434 => x"13050500",
         435 => x"6ff05fd1",
         436 => x"b7870020",
         437 => x"93870700",
         438 => x"13070040",
         439 => x"b387e740",
         440 => x"e364f5fe",
         441 => x"ef109049",
         442 => x"9307c000",
         443 => x"2320f500",
         444 => x"1305f0ff",
         445 => x"13050500",
         446 => x"6ff09fce",
         447 => x"13030500",
         448 => x"138e0500",
         449 => x"93080000",
         450 => x"63dc0500",
         451 => x"b337a000",
         452 => x"330eb040",
         453 => x"330efe40",
         454 => x"3303a040",
         455 => x"9308f0ff",
         456 => x"63dc0600",
         457 => x"b337c000",
         458 => x"b306d040",
         459 => x"93c8f8ff",
         460 => x"b386f640",
         461 => x"3306c040",
         462 => x"13070600",
         463 => x"13080300",
         464 => x"93070e00",
         465 => x"639c0628",
         466 => x"b7450000",
         467 => x"9385c598",
         468 => x"6376ce0e",
         469 => x"b7060100",
         470 => x"6378d60c",
         471 => x"93360610",
         472 => x"93b61600",
         473 => x"93963600",
         474 => x"3355d600",
         475 => x"b385a500",
         476 => x"83c50500",
         477 => x"13050002",
         478 => x"b386d500",
         479 => x"b305d540",
         480 => x"630cd500",
         481 => x"b317be00",
         482 => x"b356d300",
         483 => x"3317b600",
         484 => x"b3e7f600",
         485 => x"3318b300",
         486 => x"93550701",
         487 => x"33deb702",
         488 => x"13160701",
         489 => x"13560601",
         490 => x"b3f7b702",
         491 => x"13050e00",
         492 => x"3303c603",
         493 => x"93960701",
         494 => x"93570801",
         495 => x"b3e7d700",
         496 => x"63fe6700",
         497 => x"b307f700",
         498 => x"1305feff",
         499 => x"63e8e700",
         500 => x"63f66700",
         501 => x"1305eeff",
         502 => x"b387e700",
         503 => x"b3876740",
         504 => x"33d3b702",
         505 => x"13180801",
         506 => x"13580801",
         507 => x"b3f7b702",
         508 => x"b3066602",
         509 => x"93970701",
         510 => x"3368f800",
         511 => x"93070300",
         512 => x"637cd800",
         513 => x"33080701",
         514 => x"9307f3ff",
         515 => x"6366e800",
         516 => x"6374d800",
         517 => x"9307e3ff",
         518 => x"13150501",
         519 => x"3365f500",
         520 => x"93050000",
         521 => x"6f00000e",
         522 => x"37050001",
         523 => x"93068001",
         524 => x"e37ca6f2",
         525 => x"93060001",
         526 => x"6ff01ff3",
         527 => x"93060000",
         528 => x"630c0600",
         529 => x"b7070100",
         530 => x"637af60c",
         531 => x"93360610",
         532 => x"93b61600",
         533 => x"93963600",
         534 => x"b357d600",
         535 => x"b385f500",
         536 => x"83c70500",
         537 => x"b387d700",
         538 => x"93060002",
         539 => x"b385f640",
         540 => x"6390f60c",
         541 => x"b307ce40",
         542 => x"93051000",
         543 => x"13530701",
         544 => x"b3de6702",
         545 => x"13160701",
         546 => x"13560601",
         547 => x"93560801",
         548 => x"b3f76702",
         549 => x"13850e00",
         550 => x"330ed603",
         551 => x"93970701",
         552 => x"b3e7f600",
         553 => x"63fec701",
         554 => x"b307f700",
         555 => x"1385feff",
         556 => x"63e8e700",
         557 => x"63f6c701",
         558 => x"1385eeff",
         559 => x"b387e700",
         560 => x"b387c741",
         561 => x"33de6702",
         562 => x"13180801",
         563 => x"13580801",
         564 => x"b3f76702",
         565 => x"b306c603",
         566 => x"93970701",
         567 => x"3368f800",
         568 => x"93070e00",
         569 => x"637cd800",
         570 => x"33080701",
         571 => x"9307feff",
         572 => x"6366e800",
         573 => x"6374d800",
         574 => x"9307eeff",
         575 => x"13150501",
         576 => x"3365f500",
         577 => x"638a0800",
         578 => x"b337a000",
         579 => x"b305b040",
         580 => x"b385f540",
         581 => x"3305a040",
         582 => x"67800000",
         583 => x"b7070001",
         584 => x"93068001",
         585 => x"e37af6f2",
         586 => x"93060001",
         587 => x"6ff0dff2",
         588 => x"3317b600",
         589 => x"b356fe00",
         590 => x"13550701",
         591 => x"331ebe00",
         592 => x"b357f300",
         593 => x"b3e7c701",
         594 => x"33dea602",
         595 => x"13160701",
         596 => x"13560601",
         597 => x"3318b300",
         598 => x"b3f6a602",
         599 => x"3303c603",
         600 => x"93950601",
         601 => x"93d60701",
         602 => x"b3e6b600",
         603 => x"93050e00",
         604 => x"63fe6600",
         605 => x"b306d700",
         606 => x"9305feff",
         607 => x"63e8e600",
         608 => x"63f66600",
         609 => x"9305eeff",
         610 => x"b386e600",
         611 => x"b3866640",
         612 => x"33d3a602",
         613 => x"93970701",
         614 => x"93d70701",
         615 => x"b3f6a602",
         616 => x"33066602",
         617 => x"93960601",
         618 => x"b3e7d700",
         619 => x"93060300",
         620 => x"63fec700",
         621 => x"b307f700",
         622 => x"9306f3ff",
         623 => x"63e8e700",
         624 => x"63f6c700",
         625 => x"9306e3ff",
         626 => x"b387e700",
         627 => x"93950501",
         628 => x"b387c740",
         629 => x"b3e5d500",
         630 => x"6ff05fea",
         631 => x"6366de18",
         632 => x"b7070100",
         633 => x"63f4f604",
         634 => x"13b70610",
         635 => x"13371700",
         636 => x"13173700",
         637 => x"b7470000",
         638 => x"b3d5e600",
         639 => x"9387c798",
         640 => x"b387b700",
         641 => x"83c70700",
         642 => x"b387e700",
         643 => x"13070002",
         644 => x"b305f740",
         645 => x"6316f702",
         646 => x"13051000",
         647 => x"e3e4c6ef",
         648 => x"3335c300",
         649 => x"13351500",
         650 => x"6ff0dfed",
         651 => x"b7070001",
         652 => x"13078001",
         653 => x"e3f0f6fc",
         654 => x"13070001",
         655 => x"6ff09ffb",
         656 => x"3357f600",
         657 => x"b396b600",
         658 => x"b366d700",
         659 => x"3357fe00",
         660 => x"331ebe00",
         661 => x"b357f300",
         662 => x"b3e7c701",
         663 => x"13de0601",
         664 => x"335fc703",
         665 => x"13980601",
         666 => x"13580801",
         667 => x"3316b600",
         668 => x"3377c703",
         669 => x"b30ee803",
         670 => x"13150701",
         671 => x"13d70701",
         672 => x"3367a700",
         673 => x"13050f00",
         674 => x"637ed701",
         675 => x"3387e600",
         676 => x"1305ffff",
         677 => x"6368d700",
         678 => x"6376d701",
         679 => x"1305efff",
         680 => x"3307d700",
         681 => x"3307d741",
         682 => x"b35ec703",
         683 => x"93970701",
         684 => x"93d70701",
         685 => x"3377c703",
         686 => x"3308d803",
         687 => x"13170701",
         688 => x"b3e7e700",
         689 => x"13870e00",
         690 => x"63fe0701",
         691 => x"b387f600",
         692 => x"1387feff",
         693 => x"63e8d700",
         694 => x"63f60701",
         695 => x"1387eeff",
         696 => x"b387d700",
         697 => x"13150501",
         698 => x"b70e0100",
         699 => x"3365e500",
         700 => x"9386feff",
         701 => x"3377d500",
         702 => x"b3870741",
         703 => x"b376d600",
         704 => x"13580501",
         705 => x"13560601",
         706 => x"330ed702",
         707 => x"b306d802",
         708 => x"3307c702",
         709 => x"3308c802",
         710 => x"3306d700",
         711 => x"13570e01",
         712 => x"3307c700",
         713 => x"6374d700",
         714 => x"3308d801",
         715 => x"93560701",
         716 => x"b3860601",
         717 => x"63e6d702",
         718 => x"e394d7ce",
         719 => x"b7070100",
         720 => x"9387f7ff",
         721 => x"3377f700",
         722 => x"13170701",
         723 => x"337efe00",
         724 => x"3313b300",
         725 => x"3307c701",
         726 => x"93050000",
         727 => x"e374e3da",
         728 => x"1305f5ff",
         729 => x"6ff0dfcb",
         730 => x"93050000",
         731 => x"13050000",
         732 => x"6ff05fd9",
         733 => x"93080500",
         734 => x"13830500",
         735 => x"13070600",
         736 => x"13080500",
         737 => x"93870500",
         738 => x"63920628",
         739 => x"b7450000",
         740 => x"9385c598",
         741 => x"6376c30e",
         742 => x"b7060100",
         743 => x"6378d60c",
         744 => x"93360610",
         745 => x"93b61600",
         746 => x"93963600",
         747 => x"3355d600",
         748 => x"b385a500",
         749 => x"83c50500",
         750 => x"13050002",
         751 => x"b386d500",
         752 => x"b305d540",
         753 => x"630cd500",
         754 => x"b317b300",
         755 => x"b3d6d800",
         756 => x"3317b600",
         757 => x"b3e7f600",
         758 => x"3398b800",
         759 => x"93550701",
         760 => x"33d3b702",
         761 => x"13160701",
         762 => x"13560601",
         763 => x"b3f7b702",
         764 => x"13050300",
         765 => x"b3086602",
         766 => x"93960701",
         767 => x"93570801",
         768 => x"b3e7d700",
         769 => x"63fe1701",
         770 => x"b307f700",
         771 => x"1305f3ff",
         772 => x"63e8e700",
         773 => x"63f61701",
         774 => x"1305e3ff",
         775 => x"b387e700",
         776 => x"b3871741",
         777 => x"b3d8b702",
         778 => x"13180801",
         779 => x"13580801",
         780 => x"b3f7b702",
         781 => x"b3061603",
         782 => x"93970701",
         783 => x"3368f800",
         784 => x"93870800",
         785 => x"637cd800",
         786 => x"33080701",
         787 => x"9387f8ff",
         788 => x"6366e800",
         789 => x"6374d800",
         790 => x"9387e8ff",
         791 => x"13150501",
         792 => x"3365f500",
         793 => x"93050000",
         794 => x"67800000",
         795 => x"37050001",
         796 => x"93068001",
         797 => x"e37ca6f2",
         798 => x"93060001",
         799 => x"6ff01ff3",
         800 => x"93060000",
         801 => x"630c0600",
         802 => x"b7070100",
         803 => x"6370f60c",
         804 => x"93360610",
         805 => x"93b61600",
         806 => x"93963600",
         807 => x"b357d600",
         808 => x"b385f500",
         809 => x"83c70500",
         810 => x"b387d700",
         811 => x"93060002",
         812 => x"b385f640",
         813 => x"6396f60a",
         814 => x"b307c340",
         815 => x"93051000",
         816 => x"93580701",
         817 => x"33de1703",
         818 => x"13160701",
         819 => x"13560601",
         820 => x"93560801",
         821 => x"b3f71703",
         822 => x"13050e00",
         823 => x"3303c603",
         824 => x"93970701",
         825 => x"b3e7f600",
         826 => x"63fe6700",
         827 => x"b307f700",
         828 => x"1305feff",
         829 => x"63e8e700",
         830 => x"63f66700",
         831 => x"1305eeff",
         832 => x"b387e700",
         833 => x"b3876740",
         834 => x"33d31703",
         835 => x"13180801",
         836 => x"13580801",
         837 => x"b3f71703",
         838 => x"b3066602",
         839 => x"93970701",
         840 => x"3368f800",
         841 => x"93070300",
         842 => x"637cd800",
         843 => x"33080701",
         844 => x"9307f3ff",
         845 => x"6366e800",
         846 => x"6374d800",
         847 => x"9307e3ff",
         848 => x"13150501",
         849 => x"3365f500",
         850 => x"67800000",
         851 => x"b7070001",
         852 => x"93068001",
         853 => x"e374f6f4",
         854 => x"93060001",
         855 => x"6ff01ff4",
         856 => x"3317b600",
         857 => x"b356f300",
         858 => x"13550701",
         859 => x"3313b300",
         860 => x"b3d7f800",
         861 => x"b3e76700",
         862 => x"33d3a602",
         863 => x"13160701",
         864 => x"13560601",
         865 => x"3398b800",
         866 => x"b3f6a602",
         867 => x"b3086602",
         868 => x"93950601",
         869 => x"93d60701",
         870 => x"b3e6b600",
         871 => x"93050300",
         872 => x"63fe1601",
         873 => x"b306d700",
         874 => x"9305f3ff",
         875 => x"63e8e600",
         876 => x"63f61601",
         877 => x"9305e3ff",
         878 => x"b386e600",
         879 => x"b3861641",
         880 => x"b3d8a602",
         881 => x"93970701",
         882 => x"93d70701",
         883 => x"b3f6a602",
         884 => x"33061603",
         885 => x"93960601",
         886 => x"b3e7d700",
         887 => x"93860800",
         888 => x"63fec700",
         889 => x"b307f700",
         890 => x"9386f8ff",
         891 => x"63e8e700",
         892 => x"63f6c700",
         893 => x"9386e8ff",
         894 => x"b387e700",
         895 => x"93950501",
         896 => x"b387c740",
         897 => x"b3e5d500",
         898 => x"6ff09feb",
         899 => x"63e6d518",
         900 => x"b7070100",
         901 => x"63f4f604",
         902 => x"13b70610",
         903 => x"13371700",
         904 => x"13173700",
         905 => x"b7470000",
         906 => x"b3d5e600",
         907 => x"9387c798",
         908 => x"b387b700",
         909 => x"83c70700",
         910 => x"b387e700",
         911 => x"13070002",
         912 => x"b305f740",
         913 => x"6316f702",
         914 => x"13051000",
         915 => x"e3ee66e0",
         916 => x"33b5c800",
         917 => x"13351500",
         918 => x"67800000",
         919 => x"b7070001",
         920 => x"13078001",
         921 => x"e3f0f6fc",
         922 => x"13070001",
         923 => x"6ff09ffb",
         924 => x"3357f600",
         925 => x"b396b600",
         926 => x"b366d700",
         927 => x"3357f300",
         928 => x"3313b300",
         929 => x"b3d7f800",
         930 => x"b3e76700",
         931 => x"13d30601",
         932 => x"b35e6702",
         933 => x"13980601",
         934 => x"13580801",
         935 => x"3316b600",
         936 => x"33776702",
         937 => x"330ed803",
         938 => x"13150701",
         939 => x"13d70701",
         940 => x"3367a700",
         941 => x"13850e00",
         942 => x"637ec701",
         943 => x"3387e600",
         944 => x"1385feff",
         945 => x"6368d700",
         946 => x"6376c701",
         947 => x"1385eeff",
         948 => x"3307d700",
         949 => x"3307c741",
         950 => x"335e6702",
         951 => x"93970701",
         952 => x"93d70701",
         953 => x"33776702",
         954 => x"3308c803",
         955 => x"13170701",
         956 => x"b3e7e700",
         957 => x"13070e00",
         958 => x"63fe0701",
         959 => x"b387f600",
         960 => x"1307feff",
         961 => x"63e8d700",
         962 => x"63f60701",
         963 => x"1307eeff",
         964 => x"b387d700",
         965 => x"13150501",
         966 => x"370e0100",
         967 => x"3365e500",
         968 => x"9306feff",
         969 => x"3377d500",
         970 => x"b3870741",
         971 => x"b376d600",
         972 => x"13580501",
         973 => x"13560601",
         974 => x"3303d702",
         975 => x"b306d802",
         976 => x"3307c702",
         977 => x"3308c802",
         978 => x"3306d700",
         979 => x"13570301",
         980 => x"3307c700",
         981 => x"6374d700",
         982 => x"3308c801",
         983 => x"93560701",
         984 => x"b3860601",
         985 => x"63e6d702",
         986 => x"e39ed7ce",
         987 => x"b7070100",
         988 => x"9387f7ff",
         989 => x"3377f700",
         990 => x"13170701",
         991 => x"3373f300",
         992 => x"b398b800",
         993 => x"33076700",
         994 => x"93050000",
         995 => x"e3fee8cc",
         996 => x"1305f5ff",
         997 => x"6ff01fcd",
         998 => x"93050000",
         999 => x"13050000",
        1000 => x"67800000",
        1001 => x"13080600",
        1002 => x"93070500",
        1003 => x"13870500",
        1004 => x"63960620",
        1005 => x"b7480000",
        1006 => x"9388c898",
        1007 => x"63fcc50c",
        1008 => x"b7060100",
        1009 => x"637ed60a",
        1010 => x"93360610",
        1011 => x"93b61600",
        1012 => x"93963600",
        1013 => x"3353d600",
        1014 => x"b3886800",
        1015 => x"83c80800",
        1016 => x"13030002",
        1017 => x"b386d800",
        1018 => x"b308d340",
        1019 => x"630cd300",
        1020 => x"33971501",
        1021 => x"b356d500",
        1022 => x"33181601",
        1023 => x"33e7e600",
        1024 => x"b3171501",
        1025 => x"13560801",
        1026 => x"b356c702",
        1027 => x"13150801",
        1028 => x"13550501",
        1029 => x"3377c702",
        1030 => x"b386a602",
        1031 => x"93150701",
        1032 => x"13d70701",
        1033 => x"3367b700",
        1034 => x"637ad700",
        1035 => x"3307e800",
        1036 => x"63660701",
        1037 => x"6374d700",
        1038 => x"33070701",
        1039 => x"3307d740",
        1040 => x"b356c702",
        1041 => x"3377c702",
        1042 => x"b386a602",
        1043 => x"93970701",
        1044 => x"13170701",
        1045 => x"93d70701",
        1046 => x"b3e7e700",
        1047 => x"63fad700",
        1048 => x"b307f800",
        1049 => x"63e60701",
        1050 => x"63f4d700",
        1051 => x"b3870701",
        1052 => x"b387d740",
        1053 => x"33d51701",
        1054 => x"93050000",
        1055 => x"67800000",
        1056 => x"37030001",
        1057 => x"93068001",
        1058 => x"e37666f4",
        1059 => x"93060001",
        1060 => x"6ff05ff4",
        1061 => x"93060000",
        1062 => x"630c0600",
        1063 => x"37070100",
        1064 => x"637ee606",
        1065 => x"93360610",
        1066 => x"93b61600",
        1067 => x"93963600",
        1068 => x"3357d600",
        1069 => x"b388e800",
        1070 => x"03c70800",
        1071 => x"3307d700",
        1072 => x"93060002",
        1073 => x"b388e640",
        1074 => x"6394e606",
        1075 => x"3387c540",
        1076 => x"93550801",
        1077 => x"3356b702",
        1078 => x"13150801",
        1079 => x"13550501",
        1080 => x"93d60701",
        1081 => x"3377b702",
        1082 => x"3306a602",
        1083 => x"13170701",
        1084 => x"33e7e600",
        1085 => x"637ac700",
        1086 => x"3307e800",
        1087 => x"63660701",
        1088 => x"6374c700",
        1089 => x"33070701",
        1090 => x"3307c740",
        1091 => x"b356b702",
        1092 => x"3377b702",
        1093 => x"b386a602",
        1094 => x"6ff05ff3",
        1095 => x"37070001",
        1096 => x"93068001",
        1097 => x"e376e6f8",
        1098 => x"93060001",
        1099 => x"6ff05ff8",
        1100 => x"33181601",
        1101 => x"b3d6e500",
        1102 => x"b3171501",
        1103 => x"b3951501",
        1104 => x"3357e500",
        1105 => x"13550801",
        1106 => x"3367b700",
        1107 => x"b3d5a602",
        1108 => x"13130801",
        1109 => x"13530301",
        1110 => x"b3f6a602",
        1111 => x"b3856502",
        1112 => x"13960601",
        1113 => x"93560701",
        1114 => x"b3e6c600",
        1115 => x"63fab600",
        1116 => x"b306d800",
        1117 => x"63e60601",
        1118 => x"63f4b600",
        1119 => x"b3860601",
        1120 => x"b386b640",
        1121 => x"33d6a602",
        1122 => x"13170701",
        1123 => x"13570701",
        1124 => x"b3f6a602",
        1125 => x"33066602",
        1126 => x"93960601",
        1127 => x"3367d700",
        1128 => x"637ac700",
        1129 => x"3307e800",
        1130 => x"63660701",
        1131 => x"6374c700",
        1132 => x"33070701",
        1133 => x"3307c740",
        1134 => x"6ff09ff1",
        1135 => x"63e4d51c",
        1136 => x"37080100",
        1137 => x"63fe0605",
        1138 => x"13b80610",
        1139 => x"13381800",
        1140 => x"13183800",
        1141 => x"b7480000",
        1142 => x"33d30601",
        1143 => x"9388c898",
        1144 => x"b3886800",
        1145 => x"83c80800",
        1146 => x"13030002",
        1147 => x"b3880801",
        1148 => x"33081341",
        1149 => x"63101305",
        1150 => x"63e4b600",
        1151 => x"636cc500",
        1152 => x"3306c540",
        1153 => x"b386d540",
        1154 => x"3337c500",
        1155 => x"93070600",
        1156 => x"3387e640",
        1157 => x"13850700",
        1158 => x"93050700",
        1159 => x"67800000",
        1160 => x"b7080001",
        1161 => x"13088001",
        1162 => x"e3f616fb",
        1163 => x"13080001",
        1164 => x"6ff05ffa",
        1165 => x"b3571601",
        1166 => x"b3960601",
        1167 => x"b3e6d700",
        1168 => x"33d71501",
        1169 => x"13de0601",
        1170 => x"335fc703",
        1171 => x"13930601",
        1172 => x"13530301",
        1173 => x"b3970501",
        1174 => x"b3551501",
        1175 => x"b3e5f500",
        1176 => x"93d70501",
        1177 => x"33160601",
        1178 => x"33150501",
        1179 => x"3377c703",
        1180 => x"b30ee303",
        1181 => x"13170701",
        1182 => x"b3e7e700",
        1183 => x"13070f00",
        1184 => x"63fed701",
        1185 => x"b387f600",
        1186 => x"1307ffff",
        1187 => x"63e8d700",
        1188 => x"63f6d701",
        1189 => x"1307efff",
        1190 => x"b387d700",
        1191 => x"b387d741",
        1192 => x"b3dec703",
        1193 => x"93950501",
        1194 => x"93d50501",
        1195 => x"b3f7c703",
        1196 => x"138e0e00",
        1197 => x"3303d303",
        1198 => x"93970701",
        1199 => x"b3e5f500",
        1200 => x"63fe6500",
        1201 => x"b385b600",
        1202 => x"138efeff",
        1203 => x"63e8d500",
        1204 => x"63f66500",
        1205 => x"138eeeff",
        1206 => x"b385d500",
        1207 => x"93170701",
        1208 => x"370f0100",
        1209 => x"b3e7c701",
        1210 => x"b3856540",
        1211 => x"1303ffff",
        1212 => x"33f76700",
        1213 => x"135e0601",
        1214 => x"93d70701",
        1215 => x"33736600",
        1216 => x"b30e6702",
        1217 => x"33836702",
        1218 => x"3307c703",
        1219 => x"b387c703",
        1220 => x"330e6700",
        1221 => x"13d70e01",
        1222 => x"3307c701",
        1223 => x"63746700",
        1224 => x"b387e701",
        1225 => x"13530701",
        1226 => x"b307f300",
        1227 => x"37030100",
        1228 => x"1303f3ff",
        1229 => x"33776700",
        1230 => x"13170701",
        1231 => x"b3fe6e00",
        1232 => x"3307d701",
        1233 => x"63e6f500",
        1234 => x"639ef500",
        1235 => x"637ce500",
        1236 => x"3306c740",
        1237 => x"3333c700",
        1238 => x"b306d300",
        1239 => x"13070600",
        1240 => x"b387d740",
        1241 => x"3307e540",
        1242 => x"3335e500",
        1243 => x"b385f540",
        1244 => x"b385a540",
        1245 => x"b3981501",
        1246 => x"33570701",
        1247 => x"33e5e800",
        1248 => x"b3d50501",
        1249 => x"67800000",
        1250 => x"13030500",
        1251 => x"630a0600",
        1252 => x"2300b300",
        1253 => x"1306f6ff",
        1254 => x"13031300",
        1255 => x"e31a06fe",
        1256 => x"67800000",
        1257 => x"13030500",
        1258 => x"630e0600",
        1259 => x"83830500",
        1260 => x"23007300",
        1261 => x"1306f6ff",
        1262 => x"13031300",
        1263 => x"93851500",
        1264 => x"e31606fe",
        1265 => x"67800000",
        1266 => x"630c0602",
        1267 => x"13030500",
        1268 => x"93061000",
        1269 => x"636ab500",
        1270 => x"9306f0ff",
        1271 => x"1307f6ff",
        1272 => x"3303e300",
        1273 => x"b385e500",
        1274 => x"83830500",
        1275 => x"23007300",
        1276 => x"1306f6ff",
        1277 => x"3303d300",
        1278 => x"b385d500",
        1279 => x"e31606fe",
        1280 => x"67800000",
        1281 => x"6f000000",
        1282 => x"130101ff",
        1283 => x"23248100",
        1284 => x"13040000",
        1285 => x"23229100",
        1286 => x"23202101",
        1287 => x"23261100",
        1288 => x"93040500",
        1289 => x"13090400",
        1290 => x"93070400",
        1291 => x"732410c8",
        1292 => x"732910c0",
        1293 => x"f32710c8",
        1294 => x"e31af4fe",
        1295 => x"37460f00",
        1296 => x"13060624",
        1297 => x"93060000",
        1298 => x"13050900",
        1299 => x"93050400",
        1300 => x"eff05fb5",
        1301 => x"37460f00",
        1302 => x"23a4a400",
        1303 => x"93050400",
        1304 => x"13050900",
        1305 => x"13060624",
        1306 => x"93060000",
        1307 => x"eff08ff0",
        1308 => x"8320c100",
        1309 => x"03248100",
        1310 => x"23a0a400",
        1311 => x"23a2b400",
        1312 => x"03290100",
        1313 => x"83244100",
        1314 => x"13050000",
        1315 => x"13010101",
        1316 => x"67800000",
        1317 => x"13050000",
        1318 => x"67800000",
        1319 => x"13050000",
        1320 => x"67800000",
        1321 => x"130101ff",
        1322 => x"23202101",
        1323 => x"23261100",
        1324 => x"13090600",
        1325 => x"6356c002",
        1326 => x"23248100",
        1327 => x"23229100",
        1328 => x"13840500",
        1329 => x"b384c500",
        1330 => x"03450400",
        1331 => x"13041400",
        1332 => x"efe0dfba",
        1333 => x"e39a84fe",
        1334 => x"03248100",
        1335 => x"83244100",
        1336 => x"8320c100",
        1337 => x"13050900",
        1338 => x"03290100",
        1339 => x"13010101",
        1340 => x"67800000",
        1341 => x"130101ff",
        1342 => x"23202101",
        1343 => x"23261100",
        1344 => x"13090600",
        1345 => x"6356c002",
        1346 => x"23248100",
        1347 => x"23229100",
        1348 => x"13840500",
        1349 => x"b384c500",
        1350 => x"efe01fb6",
        1351 => x"13041400",
        1352 => x"a30fa4fe",
        1353 => x"e39a84fe",
        1354 => x"03248100",
        1355 => x"83244100",
        1356 => x"8320c100",
        1357 => x"13050900",
        1358 => x"03290100",
        1359 => x"13010101",
        1360 => x"67800000",
        1361 => x"13051000",
        1362 => x"67800000",
        1363 => x"130101ff",
        1364 => x"23261100",
        1365 => x"ef009062",
        1366 => x"8320c100",
        1367 => x"93076001",
        1368 => x"2320f500",
        1369 => x"1305f0ff",
        1370 => x"13010101",
        1371 => x"67800000",
        1372 => x"1305f0ff",
        1373 => x"67800000",
        1374 => x"b7270000",
        1375 => x"23a2f500",
        1376 => x"13050000",
        1377 => x"67800000",
        1378 => x"13051000",
        1379 => x"67800000",
        1380 => x"13050000",
        1381 => x"67800000",
        1382 => x"130101fe",
        1383 => x"2324c100",
        1384 => x"2326d100",
        1385 => x"2328e100",
        1386 => x"232af100",
        1387 => x"232c0101",
        1388 => x"232e1101",
        1389 => x"1305f0ff",
        1390 => x"13010102",
        1391 => x"67800000",
        1392 => x"130101ff",
        1393 => x"23261100",
        1394 => x"ef00505b",
        1395 => x"8320c100",
        1396 => x"9307a000",
        1397 => x"2320f500",
        1398 => x"1305f0ff",
        1399 => x"13010101",
        1400 => x"67800000",
        1401 => x"130101ff",
        1402 => x"23261100",
        1403 => x"ef001059",
        1404 => x"8320c100",
        1405 => x"93072000",
        1406 => x"2320f500",
        1407 => x"1305f0ff",
        1408 => x"13010101",
        1409 => x"67800000",
        1410 => x"b7270000",
        1411 => x"23a2f500",
        1412 => x"13050000",
        1413 => x"67800000",
        1414 => x"130101ff",
        1415 => x"23261100",
        1416 => x"ef00d055",
        1417 => x"8320c100",
        1418 => x"9307f001",
        1419 => x"2320f500",
        1420 => x"1305f0ff",
        1421 => x"13010101",
        1422 => x"67800000",
        1423 => x"130101ff",
        1424 => x"23261100",
        1425 => x"ef009053",
        1426 => x"8320c100",
        1427 => x"9307b000",
        1428 => x"2320f500",
        1429 => x"1305f0ff",
        1430 => x"13010101",
        1431 => x"67800000",
        1432 => x"130101ff",
        1433 => x"23261100",
        1434 => x"ef005051",
        1435 => x"8320c100",
        1436 => x"9307c000",
        1437 => x"2320f500",
        1438 => x"1305f0ff",
        1439 => x"13010101",
        1440 => x"67800000",
        1441 => x"03a7c187",
        1442 => x"b7870020",
        1443 => x"93870700",
        1444 => x"93060040",
        1445 => x"b387d740",
        1446 => x"630c0700",
        1447 => x"3305a700",
        1448 => x"63e2a702",
        1449 => x"23aea186",
        1450 => x"13050700",
        1451 => x"67800000",
        1452 => x"9386819c",
        1453 => x"1387819c",
        1454 => x"23aed186",
        1455 => x"3305a700",
        1456 => x"e3f2a7fe",
        1457 => x"130101ff",
        1458 => x"23261100",
        1459 => x"ef00104b",
        1460 => x"8320c100",
        1461 => x"9307c000",
        1462 => x"2320f500",
        1463 => x"1307f0ff",
        1464 => x"13050700",
        1465 => x"13010101",
        1466 => x"67800000",
        1467 => x"370700f0",
        1468 => x"13070702",
        1469 => x"83274700",
        1470 => x"93f74700",
        1471 => x"e38c07fe",
        1472 => x"03258700",
        1473 => x"1375f50f",
        1474 => x"67800000",
        1475 => x"f32710fc",
        1476 => x"63960700",
        1477 => x"b7f7fa02",
        1478 => x"93870708",
        1479 => x"63060500",
        1480 => x"33d5a702",
        1481 => x"1305f5ff",
        1482 => x"b70700f0",
        1483 => x"23a6a702",
        1484 => x"23a0b702",
        1485 => x"67800000",
        1486 => x"370700f0",
        1487 => x"1375f50f",
        1488 => x"13070702",
        1489 => x"2324a700",
        1490 => x"83274700",
        1491 => x"93f70701",
        1492 => x"e38c07fe",
        1493 => x"67800000",
        1494 => x"630e0502",
        1495 => x"130101ff",
        1496 => x"23248100",
        1497 => x"23261100",
        1498 => x"13040500",
        1499 => x"03450500",
        1500 => x"630a0500",
        1501 => x"13041400",
        1502 => x"eff01ffc",
        1503 => x"03450400",
        1504 => x"e31a05fe",
        1505 => x"8320c100",
        1506 => x"03248100",
        1507 => x"13010101",
        1508 => x"67800000",
        1509 => x"67800000",
        1510 => x"130101f9",
        1511 => x"23229106",
        1512 => x"23202107",
        1513 => x"23261106",
        1514 => x"23248106",
        1515 => x"232e3105",
        1516 => x"232c4105",
        1517 => x"232a5105",
        1518 => x"23286105",
        1519 => x"23267105",
        1520 => x"23248105",
        1521 => x"23229105",
        1522 => x"2320a105",
        1523 => x"13090500",
        1524 => x"93840500",
        1525 => x"232c0100",
        1526 => x"232e0100",
        1527 => x"23200102",
        1528 => x"23220102",
        1529 => x"23240102",
        1530 => x"23260102",
        1531 => x"23280102",
        1532 => x"232a0102",
        1533 => x"232c0102",
        1534 => x"232e0102",
        1535 => x"732410fc",
        1536 => x"63160400",
        1537 => x"37f4fa02",
        1538 => x"13040408",
        1539 => x"97f2ffff",
        1540 => x"938282af",
        1541 => x"73905230",
        1542 => x"37c50100",
        1543 => x"93050004",
        1544 => x"13050520",
        1545 => x"eff09fee",
        1546 => x"b7270000",
        1547 => x"93870771",
        1548 => x"b356f402",
        1549 => x"13561400",
        1550 => x"370700f0",
        1551 => x"1306f6ff",
        1552 => x"b7170300",
        1553 => x"2326c708",
        1554 => x"130e1001",
        1555 => x"938707d4",
        1556 => x"2320c709",
        1557 => x"370600f0",
        1558 => x"37230000",
        1559 => x"1303f370",
        1560 => x"37581200",
        1561 => x"130808f8",
        1562 => x"b70800f0",
        1563 => x"370500f0",
        1564 => x"b70500f0",
        1565 => x"3357f402",
        1566 => x"9387f6ff",
        1567 => x"2328f60a",
        1568 => x"2326660a",
        1569 => x"2320c60b",
        1570 => x"93078070",
        1571 => x"23a0f806",
        1572 => x"b3570403",
        1573 => x"1307f7ff",
        1574 => x"13170701",
        1575 => x"13678700",
        1576 => x"2320e504",
        1577 => x"1307a007",
        1578 => x"9387f7ff",
        1579 => x"93970701",
        1580 => x"93e7c700",
        1581 => x"23a8f504",
        1582 => x"b70700f0",
        1583 => x"23ace700",
        1584 => x"f3224030",
        1585 => x"93e20208",
        1586 => x"73904230",
        1587 => x"f3224030",
        1588 => x"93e28200",
        1589 => x"73904230",
        1590 => x"b7220000",
        1591 => x"93828280",
        1592 => x"73900230",
        1593 => x"b7490000",
        1594 => x"1385c9aa",
        1595 => x"eff0dfe6",
        1596 => x"1304f9ff",
        1597 => x"63522003",
        1598 => x"1309f0ff",
        1599 => x"03a50400",
        1600 => x"1304f4ff",
        1601 => x"93844400",
        1602 => x"eff01fe5",
        1603 => x"1385c9aa",
        1604 => x"eff09fe4",
        1605 => x"e31424ff",
        1606 => x"37450000",
        1607 => x"130505ab",
        1608 => x"37f9eeee",
        1609 => x"b7faeeee",
        1610 => x"b7090010",
        1611 => x"37140000",
        1612 => x"eff09fe2",
        1613 => x"374b0000",
        1614 => x"9389f9ff",
        1615 => x"1309f9ee",
        1616 => x"938aeaee",
        1617 => x"130404e1",
        1618 => x"93040000",
        1619 => x"b71b0000",
        1620 => x"938b0b2c",
        1621 => x"130af000",
        1622 => x"6f00c000",
        1623 => x"938bfbff",
        1624 => x"63840b18",
        1625 => x"93050000",
        1626 => x"13058100",
        1627 => x"ef00502b",
        1628 => x"e31605fe",
        1629 => x"032c8100",
        1630 => x"8325c100",
        1631 => x"13060400",
        1632 => x"9357cc01",
        1633 => x"13974500",
        1634 => x"b367f700",
        1635 => x"b3f73701",
        1636 => x"33773c01",
        1637 => x"13d5f541",
        1638 => x"13d88501",
        1639 => x"3307f700",
        1640 => x"33070701",
        1641 => x"9377d500",
        1642 => x"3307f700",
        1643 => x"33774703",
        1644 => x"937725ff",
        1645 => x"93860400",
        1646 => x"13050c00",
        1647 => x"938bfbff",
        1648 => x"3307f700",
        1649 => x"b307ec40",
        1650 => x"1357f741",
        1651 => x"3338fc00",
        1652 => x"3387e540",
        1653 => x"33070741",
        1654 => x"b3885703",
        1655 => x"33072703",
        1656 => x"33b82703",
        1657 => x"33071701",
        1658 => x"b3872703",
        1659 => x"33070701",
        1660 => x"1358f741",
        1661 => x"13783800",
        1662 => x"b307f800",
        1663 => x"33b80701",
        1664 => x"3307e800",
        1665 => x"1318e701",
        1666 => x"93d72700",
        1667 => x"b367f800",
        1668 => x"13582740",
        1669 => x"93184800",
        1670 => x"13d3c701",
        1671 => x"33e36800",
        1672 => x"33733301",
        1673 => x"b3f83701",
        1674 => x"135e8801",
        1675 => x"1357f741",
        1676 => x"b3886800",
        1677 => x"b388c801",
        1678 => x"1373d700",
        1679 => x"b3886800",
        1680 => x"b3f84803",
        1681 => x"137727ff",
        1682 => x"939c4700",
        1683 => x"b38cfc40",
        1684 => x"939c2c00",
        1685 => x"b30c9c41",
        1686 => x"b388e800",
        1687 => x"33871741",
        1688 => x"93d8f841",
        1689 => x"33b3e700",
        1690 => x"33081841",
        1691 => x"33086840",
        1692 => x"33082803",
        1693 => x"33035703",
        1694 => x"b3382703",
        1695 => x"33086800",
        1696 => x"33072703",
        1697 => x"33081801",
        1698 => x"9358f841",
        1699 => x"93f83800",
        1700 => x"3387e800",
        1701 => x"b3381701",
        1702 => x"b3880801",
        1703 => x"9398e801",
        1704 => x"13572700",
        1705 => x"33e7e800",
        1706 => x"13184700",
        1707 => x"3307e840",
        1708 => x"13172700",
        1709 => x"338de740",
        1710 => x"efe05fc4",
        1711 => x"83260101",
        1712 => x"13070500",
        1713 => x"13880c00",
        1714 => x"93070d00",
        1715 => x"13060c00",
        1716 => x"93050bae",
        1717 => x"13058101",
        1718 => x"ef008046",
        1719 => x"13058101",
        1720 => x"eff09fc7",
        1721 => x"e3900be8",
        1722 => x"73001000",
        1723 => x"b70700f0",
        1724 => x"9306f00f",
        1725 => x"23a4d706",
        1726 => x"370700f0",
        1727 => x"83260704",
        1728 => x"93050009",
        1729 => x"b70700f0",
        1730 => x"93e60630",
        1731 => x"2320d704",
        1732 => x"2324b704",
        1733 => x"03a60705",
        1734 => x"b70600f0",
        1735 => x"13660630",
        1736 => x"23a8c704",
        1737 => x"23acb704",
        1738 => x"93071000",
        1739 => x"23a6f60e",
        1740 => x"6ff0dfe1",
        1741 => x"130101ff",
        1742 => x"23248100",
        1743 => x"23261100",
        1744 => x"93070000",
        1745 => x"13040500",
        1746 => x"63880700",
        1747 => x"93050000",
        1748 => x"97000000",
        1749 => x"e7000000",
        1750 => x"83a70188",
        1751 => x"63840700",
        1752 => x"e7800700",
        1753 => x"13050400",
        1754 => x"eff0df89",
        1755 => x"13050000",
        1756 => x"67800000",
        1757 => x"130101ff",
        1758 => x"23248100",
        1759 => x"23261100",
        1760 => x"13040500",
        1761 => x"2316b500",
        1762 => x"2317c500",
        1763 => x"23200500",
        1764 => x"23220500",
        1765 => x"23240500",
        1766 => x"23220506",
        1767 => x"23280500",
        1768 => x"232a0500",
        1769 => x"232c0500",
        1770 => x"13068000",
        1771 => x"93050000",
        1772 => x"1305c505",
        1773 => x"eff04ffd",
        1774 => x"b7270000",
        1775 => x"938707fb",
        1776 => x"2322f402",
        1777 => x"b7270000",
        1778 => x"93878700",
        1779 => x"2324f402",
        1780 => x"b7270000",
        1781 => x"9387c708",
        1782 => x"2326f402",
        1783 => x"b7270000",
        1784 => x"9387470e",
        1785 => x"8320c100",
        1786 => x"23208402",
        1787 => x"2328f402",
        1788 => x"03248100",
        1789 => x"13010101",
        1790 => x"67800000",
        1791 => x"b7350000",
        1792 => x"37050020",
        1793 => x"13868181",
        1794 => x"9385c555",
        1795 => x"13054502",
        1796 => x"6f00c021",
        1797 => x"83254500",
        1798 => x"130101ff",
        1799 => x"b7070020",
        1800 => x"23248100",
        1801 => x"23261100",
        1802 => x"93870709",
        1803 => x"13040500",
        1804 => x"6384f500",
        1805 => x"ef109012",
        1806 => x"83258400",
        1807 => x"9387818f",
        1808 => x"6386f500",
        1809 => x"13050400",
        1810 => x"ef105011",
        1811 => x"8325c400",
        1812 => x"93870196",
        1813 => x"638cf500",
        1814 => x"13050400",
        1815 => x"03248100",
        1816 => x"8320c100",
        1817 => x"13010101",
        1818 => x"6f10500f",
        1819 => x"8320c100",
        1820 => x"03248100",
        1821 => x"13010101",
        1822 => x"67800000",
        1823 => x"b7270000",
        1824 => x"37050020",
        1825 => x"130101ff",
        1826 => x"9387c7bf",
        1827 => x"13060000",
        1828 => x"93054000",
        1829 => x"13050509",
        1830 => x"23261100",
        1831 => x"23a0f188",
        1832 => x"eff05fed",
        1833 => x"13061000",
        1834 => x"93059000",
        1835 => x"1385818f",
        1836 => x"eff05fec",
        1837 => x"8320c100",
        1838 => x"13062000",
        1839 => x"93052001",
        1840 => x"13850196",
        1841 => x"13010101",
        1842 => x"6ff0dfea",
        1843 => x"13050000",
        1844 => x"67800000",
        1845 => x"83a70188",
        1846 => x"130101ff",
        1847 => x"23202101",
        1848 => x"23261100",
        1849 => x"23248100",
        1850 => x"23229100",
        1851 => x"13090500",
        1852 => x"63940700",
        1853 => x"eff09ff8",
        1854 => x"93848181",
        1855 => x"03a48400",
        1856 => x"83a74400",
        1857 => x"9387f7ff",
        1858 => x"63d80702",
        1859 => x"83a70400",
        1860 => x"6390070c",
        1861 => x"9305c01a",
        1862 => x"13050900",
        1863 => x"ef001009",
        1864 => x"13040500",
        1865 => x"63140508",
        1866 => x"23a00400",
        1867 => x"9307c000",
        1868 => x"2320f900",
        1869 => x"6f004005",
        1870 => x"0317c400",
        1871 => x"63140706",
        1872 => x"b707ffff",
        1873 => x"93871700",
        1874 => x"23220406",
        1875 => x"23200400",
        1876 => x"23220400",
        1877 => x"23240400",
        1878 => x"2326f400",
        1879 => x"23280400",
        1880 => x"232a0400",
        1881 => x"232c0400",
        1882 => x"13068000",
        1883 => x"93050000",
        1884 => x"1305c405",
        1885 => x"eff04fe1",
        1886 => x"232a0402",
        1887 => x"232c0402",
        1888 => x"23240404",
        1889 => x"23260404",
        1890 => x"8320c100",
        1891 => x"13050400",
        1892 => x"03248100",
        1893 => x"83244100",
        1894 => x"03290100",
        1895 => x"13010101",
        1896 => x"67800000",
        1897 => x"13048406",
        1898 => x"6ff0dff5",
        1899 => x"93074000",
        1900 => x"23200500",
        1901 => x"2322f500",
        1902 => x"1305c500",
        1903 => x"2324a400",
        1904 => x"1306001a",
        1905 => x"93050000",
        1906 => x"eff00fdc",
        1907 => x"23a08400",
        1908 => x"83a40400",
        1909 => x"6ff09ff2",
        1910 => x"83270502",
        1911 => x"639e0700",
        1912 => x"b7270000",
        1913 => x"938747c1",
        1914 => x"2320f502",
        1915 => x"83a70188",
        1916 => x"63940700",
        1917 => x"6ff09fe8",
        1918 => x"67800000",
        1919 => x"67800000",
        1920 => x"67800000",
        1921 => x"b7250000",
        1922 => x"13868181",
        1923 => x"9385c5b6",
        1924 => x"13050000",
        1925 => x"6f008001",
        1926 => x"b7250000",
        1927 => x"13868181",
        1928 => x"9385c5cc",
        1929 => x"13050000",
        1930 => x"6f004000",
        1931 => x"130101fd",
        1932 => x"23248102",
        1933 => x"23202103",
        1934 => x"232e3101",
        1935 => x"232c4101",
        1936 => x"23286101",
        1937 => x"23267101",
        1938 => x"23261102",
        1939 => x"23229102",
        1940 => x"232a5101",
        1941 => x"93090500",
        1942 => x"138a0500",
        1943 => x"13040600",
        1944 => x"13090000",
        1945 => x"130b1000",
        1946 => x"930bf0ff",
        1947 => x"83248400",
        1948 => x"832a4400",
        1949 => x"938afaff",
        1950 => x"63de0a02",
        1951 => x"03240400",
        1952 => x"e31604fe",
        1953 => x"8320c102",
        1954 => x"03248102",
        1955 => x"83244102",
        1956 => x"8329c101",
        1957 => x"032a8101",
        1958 => x"832a4101",
        1959 => x"032b0101",
        1960 => x"832bc100",
        1961 => x"13050900",
        1962 => x"03290102",
        1963 => x"13010103",
        1964 => x"67800000",
        1965 => x"83d7c400",
        1966 => x"637efb00",
        1967 => x"8397e400",
        1968 => x"638a7701",
        1969 => x"93850400",
        1970 => x"13850900",
        1971 => x"e7000a00",
        1972 => x"3369a900",
        1973 => x"93848406",
        1974 => x"6ff0dff9",
        1975 => x"130101f6",
        1976 => x"232af108",
        1977 => x"b7070080",
        1978 => x"9387f7ff",
        1979 => x"232ef100",
        1980 => x"2328f100",
        1981 => x"b707ffff",
        1982 => x"2326d108",
        1983 => x"2324b100",
        1984 => x"232cb100",
        1985 => x"93878720",
        1986 => x"9306c108",
        1987 => x"93058100",
        1988 => x"232e1106",
        1989 => x"232af100",
        1990 => x"2328e108",
        1991 => x"232c0109",
        1992 => x"232e1109",
        1993 => x"2322d100",
        1994 => x"ef00d037",
        1995 => x"83278100",
        1996 => x"23800700",
        1997 => x"8320c107",
        1998 => x"1301010a",
        1999 => x"67800000",
        2000 => x"130101f6",
        2001 => x"232af108",
        2002 => x"b7070080",
        2003 => x"9387f7ff",
        2004 => x"232ef100",
        2005 => x"2328f100",
        2006 => x"b707ffff",
        2007 => x"93878720",
        2008 => x"232af100",
        2009 => x"2324a100",
        2010 => x"232ca100",
        2011 => x"03a54187",
        2012 => x"2324c108",
        2013 => x"2326d108",
        2014 => x"13860500",
        2015 => x"93068108",
        2016 => x"93058100",
        2017 => x"232e1106",
        2018 => x"2328e108",
        2019 => x"232c0109",
        2020 => x"232e1109",
        2021 => x"2322d100",
        2022 => x"ef00d030",
        2023 => x"83278100",
        2024 => x"23800700",
        2025 => x"8320c107",
        2026 => x"1301010a",
        2027 => x"67800000",
        2028 => x"130101ff",
        2029 => x"23248100",
        2030 => x"13840500",
        2031 => x"8395e500",
        2032 => x"23261100",
        2033 => x"ef008031",
        2034 => x"63400502",
        2035 => x"83274405",
        2036 => x"b387a700",
        2037 => x"232af404",
        2038 => x"8320c100",
        2039 => x"03248100",
        2040 => x"13010101",
        2041 => x"67800000",
        2042 => x"8357c400",
        2043 => x"37f7ffff",
        2044 => x"1307f7ff",
        2045 => x"b3f7e700",
        2046 => x"2316f400",
        2047 => x"6ff0dffd",
        2048 => x"13050000",
        2049 => x"67800000",
        2050 => x"83d7c500",
        2051 => x"130101fe",
        2052 => x"232c8100",
        2053 => x"232a9100",
        2054 => x"23282101",
        2055 => x"23263101",
        2056 => x"232e1100",
        2057 => x"93f70710",
        2058 => x"93040500",
        2059 => x"13840500",
        2060 => x"13090600",
        2061 => x"93890600",
        2062 => x"638a0700",
        2063 => x"8395e500",
        2064 => x"93062000",
        2065 => x"13060000",
        2066 => x"ef004024",
        2067 => x"8357c400",
        2068 => x"37f7ffff",
        2069 => x"1307f7ff",
        2070 => x"b3f7e700",
        2071 => x"8315e400",
        2072 => x"2316f400",
        2073 => x"03248101",
        2074 => x"8320c101",
        2075 => x"93860900",
        2076 => x"13060900",
        2077 => x"8329c100",
        2078 => x"03290101",
        2079 => x"13850400",
        2080 => x"83244101",
        2081 => x"13010102",
        2082 => x"6f00402a",
        2083 => x"130101ff",
        2084 => x"23248100",
        2085 => x"13840500",
        2086 => x"8395e500",
        2087 => x"23261100",
        2088 => x"ef00c01e",
        2089 => x"1307f0ff",
        2090 => x"8357c400",
        2091 => x"6312e502",
        2092 => x"37f7ffff",
        2093 => x"1307f7ff",
        2094 => x"b3f7e700",
        2095 => x"2316f400",
        2096 => x"8320c100",
        2097 => x"03248100",
        2098 => x"13010101",
        2099 => x"67800000",
        2100 => x"37170000",
        2101 => x"b3e7e700",
        2102 => x"2316f400",
        2103 => x"232aa404",
        2104 => x"6ff01ffe",
        2105 => x"8395e500",
        2106 => x"6f004000",
        2107 => x"130101ff",
        2108 => x"23248100",
        2109 => x"23229100",
        2110 => x"13040500",
        2111 => x"13850500",
        2112 => x"23261100",
        2113 => x"23a20188",
        2114 => x"eff08fc6",
        2115 => x"9307f0ff",
        2116 => x"6318f500",
        2117 => x"83a74188",
        2118 => x"63840700",
        2119 => x"2320f400",
        2120 => x"8320c100",
        2121 => x"03248100",
        2122 => x"83244100",
        2123 => x"13010101",
        2124 => x"67800000",
        2125 => x"83a74187",
        2126 => x"6388a714",
        2127 => x"8327c501",
        2128 => x"130101fe",
        2129 => x"232c8100",
        2130 => x"232e1100",
        2131 => x"232a9100",
        2132 => x"23282101",
        2133 => x"23263101",
        2134 => x"13040500",
        2135 => x"638a0704",
        2136 => x"83a7c700",
        2137 => x"638c0702",
        2138 => x"93040000",
        2139 => x"13090008",
        2140 => x"8327c401",
        2141 => x"83a7c700",
        2142 => x"b3879700",
        2143 => x"83a50700",
        2144 => x"639c050c",
        2145 => x"93844400",
        2146 => x"e39424ff",
        2147 => x"8327c401",
        2148 => x"13050400",
        2149 => x"83a5c700",
        2150 => x"ef008029",
        2151 => x"8327c401",
        2152 => x"83a50700",
        2153 => x"63860500",
        2154 => x"13050400",
        2155 => x"ef004028",
        2156 => x"83254401",
        2157 => x"63860500",
        2158 => x"13050400",
        2159 => x"ef004027",
        2160 => x"8325c401",
        2161 => x"63860500",
        2162 => x"13050400",
        2163 => x"ef004026",
        2164 => x"83250403",
        2165 => x"63860500",
        2166 => x"13050400",
        2167 => x"ef004025",
        2168 => x"83254403",
        2169 => x"63860500",
        2170 => x"13050400",
        2171 => x"ef004024",
        2172 => x"83258403",
        2173 => x"63860500",
        2174 => x"13050400",
        2175 => x"ef004023",
        2176 => x"83258404",
        2177 => x"63860500",
        2178 => x"13050400",
        2179 => x"ef004022",
        2180 => x"83254404",
        2181 => x"63860500",
        2182 => x"13050400",
        2183 => x"ef004021",
        2184 => x"8325c402",
        2185 => x"63860500",
        2186 => x"13050400",
        2187 => x"ef004020",
        2188 => x"83270402",
        2189 => x"638c0702",
        2190 => x"13050400",
        2191 => x"03248101",
        2192 => x"8320c101",
        2193 => x"83244101",
        2194 => x"03290101",
        2195 => x"8329c100",
        2196 => x"13010102",
        2197 => x"67800700",
        2198 => x"83a90500",
        2199 => x"13050400",
        2200 => x"ef00001d",
        2201 => x"93850900",
        2202 => x"6ff09ff1",
        2203 => x"8320c101",
        2204 => x"03248101",
        2205 => x"83244101",
        2206 => x"03290101",
        2207 => x"8329c100",
        2208 => x"13010102",
        2209 => x"67800000",
        2210 => x"67800000",
        2211 => x"130101ff",
        2212 => x"23248100",
        2213 => x"23229100",
        2214 => x"13040500",
        2215 => x"13850500",
        2216 => x"93050600",
        2217 => x"13860600",
        2218 => x"23261100",
        2219 => x"23a20188",
        2220 => x"eff00fae",
        2221 => x"9307f0ff",
        2222 => x"6318f500",
        2223 => x"83a74188",
        2224 => x"63840700",
        2225 => x"2320f400",
        2226 => x"8320c100",
        2227 => x"03248100",
        2228 => x"83244100",
        2229 => x"13010101",
        2230 => x"67800000",
        2231 => x"130101ff",
        2232 => x"23248100",
        2233 => x"23229100",
        2234 => x"13040500",
        2235 => x"13850500",
        2236 => x"93050600",
        2237 => x"13860600",
        2238 => x"23261100",
        2239 => x"23a20188",
        2240 => x"eff04f9f",
        2241 => x"9307f0ff",
        2242 => x"6318f500",
        2243 => x"83a74188",
        2244 => x"63840700",
        2245 => x"2320f400",
        2246 => x"8320c100",
        2247 => x"03248100",
        2248 => x"83244100",
        2249 => x"13010101",
        2250 => x"67800000",
        2251 => x"130101ff",
        2252 => x"23248100",
        2253 => x"23229100",
        2254 => x"13040500",
        2255 => x"13850500",
        2256 => x"93050600",
        2257 => x"13860600",
        2258 => x"23261100",
        2259 => x"23a20188",
        2260 => x"eff04f95",
        2261 => x"9307f0ff",
        2262 => x"6318f500",
        2263 => x"83a74188",
        2264 => x"63840700",
        2265 => x"2320f400",
        2266 => x"8320c100",
        2267 => x"03248100",
        2268 => x"83244100",
        2269 => x"13010101",
        2270 => x"67800000",
        2271 => x"03a54187",
        2272 => x"67800000",
        2273 => x"130101ff",
        2274 => x"23248100",
        2275 => x"23229100",
        2276 => x"37440000",
        2277 => x"b7440000",
        2278 => x"938704c4",
        2279 => x"130404c4",
        2280 => x"3304f440",
        2281 => x"23202101",
        2282 => x"23261100",
        2283 => x"13542440",
        2284 => x"938404c4",
        2285 => x"13090000",
        2286 => x"63108904",
        2287 => x"b7440000",
        2288 => x"37440000",
        2289 => x"938704c4",
        2290 => x"130404c4",
        2291 => x"3304f440",
        2292 => x"13542440",
        2293 => x"938404c4",
        2294 => x"13090000",
        2295 => x"63188902",
        2296 => x"8320c100",
        2297 => x"03248100",
        2298 => x"83244100",
        2299 => x"03290100",
        2300 => x"13010101",
        2301 => x"67800000",
        2302 => x"83a70400",
        2303 => x"13091900",
        2304 => x"93844400",
        2305 => x"e7800700",
        2306 => x"6ff01ffb",
        2307 => x"83a70400",
        2308 => x"13091900",
        2309 => x"93844400",
        2310 => x"e7800700",
        2311 => x"6ff01ffc",
        2312 => x"13860500",
        2313 => x"93050500",
        2314 => x"03a54187",
        2315 => x"6f10401e",
        2316 => x"638a050e",
        2317 => x"83a7c5ff",
        2318 => x"130101fe",
        2319 => x"232c8100",
        2320 => x"232e1100",
        2321 => x"1384c5ff",
        2322 => x"63d40700",
        2323 => x"3304f400",
        2324 => x"2326a100",
        2325 => x"ef008031",
        2326 => x"83a7c188",
        2327 => x"0325c100",
        2328 => x"639e0700",
        2329 => x"23220400",
        2330 => x"23a68188",
        2331 => x"03248101",
        2332 => x"8320c101",
        2333 => x"13010102",
        2334 => x"6f00802f",
        2335 => x"6374f402",
        2336 => x"03260400",
        2337 => x"b306c400",
        2338 => x"639ad700",
        2339 => x"83a60700",
        2340 => x"83a74700",
        2341 => x"b386c600",
        2342 => x"2320d400",
        2343 => x"2322f400",
        2344 => x"6ff09ffc",
        2345 => x"13870700",
        2346 => x"83a74700",
        2347 => x"63840700",
        2348 => x"e37af4fe",
        2349 => x"83260700",
        2350 => x"3306d700",
        2351 => x"63188602",
        2352 => x"03260400",
        2353 => x"b386c600",
        2354 => x"2320d700",
        2355 => x"3306d700",
        2356 => x"e39ec7f8",
        2357 => x"03a60700",
        2358 => x"83a74700",
        2359 => x"b306d600",
        2360 => x"2320d700",
        2361 => x"2322f700",
        2362 => x"6ff05ff8",
        2363 => x"6378c400",
        2364 => x"9307c000",
        2365 => x"2320f500",
        2366 => x"6ff05ff7",
        2367 => x"03260400",
        2368 => x"b306c400",
        2369 => x"639ad700",
        2370 => x"83a60700",
        2371 => x"83a74700",
        2372 => x"b386c600",
        2373 => x"2320d400",
        2374 => x"2322f400",
        2375 => x"23228700",
        2376 => x"6ff0dff4",
        2377 => x"67800000",
        2378 => x"130101ff",
        2379 => x"23202101",
        2380 => x"83a78188",
        2381 => x"23248100",
        2382 => x"23229100",
        2383 => x"23261100",
        2384 => x"93040500",
        2385 => x"13840500",
        2386 => x"63980700",
        2387 => x"93050000",
        2388 => x"ef10c010",
        2389 => x"23a4a188",
        2390 => x"93050400",
        2391 => x"13850400",
        2392 => x"ef10c00f",
        2393 => x"1309f0ff",
        2394 => x"63122503",
        2395 => x"1304f0ff",
        2396 => x"8320c100",
        2397 => x"13050400",
        2398 => x"03248100",
        2399 => x"83244100",
        2400 => x"03290100",
        2401 => x"13010101",
        2402 => x"67800000",
        2403 => x"13043500",
        2404 => x"1374c4ff",
        2405 => x"e30e85fc",
        2406 => x"b305a440",
        2407 => x"13850400",
        2408 => x"ef10c00b",
        2409 => x"e31625fd",
        2410 => x"6ff05ffc",
        2411 => x"130101fe",
        2412 => x"232a9100",
        2413 => x"93843500",
        2414 => x"93f4c4ff",
        2415 => x"23282101",
        2416 => x"232e1100",
        2417 => x"232c8100",
        2418 => x"23263101",
        2419 => x"23244101",
        2420 => x"93848400",
        2421 => x"9307c000",
        2422 => x"13090500",
        2423 => x"63f0f40a",
        2424 => x"9304c000",
        2425 => x"63eeb408",
        2426 => x"13050900",
        2427 => x"ef000018",
        2428 => x"83a7c188",
        2429 => x"13840700",
        2430 => x"631a040a",
        2431 => x"93850400",
        2432 => x"13050900",
        2433 => x"eff05ff2",
        2434 => x"9307f0ff",
        2435 => x"13040500",
        2436 => x"6316f514",
        2437 => x"03a4c188",
        2438 => x"93070400",
        2439 => x"639c0710",
        2440 => x"63040412",
        2441 => x"032a0400",
        2442 => x"93050000",
        2443 => x"13050900",
        2444 => x"330a4401",
        2445 => x"ef108002",
        2446 => x"6318aa10",
        2447 => x"83270400",
        2448 => x"13050900",
        2449 => x"b384f440",
        2450 => x"93850400",
        2451 => x"eff0dfed",
        2452 => x"9307f0ff",
        2453 => x"630af50e",
        2454 => x"83270400",
        2455 => x"b3879700",
        2456 => x"2320f400",
        2457 => x"83a7c188",
        2458 => x"638e070e",
        2459 => x"03a74700",
        2460 => x"6318870c",
        2461 => x"23a20700",
        2462 => x"6f004006",
        2463 => x"e3d404f6",
        2464 => x"9307c000",
        2465 => x"2320f900",
        2466 => x"13050000",
        2467 => x"8320c101",
        2468 => x"03248101",
        2469 => x"83244101",
        2470 => x"03290101",
        2471 => x"8329c100",
        2472 => x"032a8100",
        2473 => x"13010102",
        2474 => x"67800000",
        2475 => x"83260400",
        2476 => x"b3869640",
        2477 => x"63ca0606",
        2478 => x"1307b000",
        2479 => x"637ad704",
        2480 => x"23209400",
        2481 => x"33079400",
        2482 => x"63908704",
        2483 => x"23a6e188",
        2484 => x"83274400",
        2485 => x"2320d700",
        2486 => x"2322f700",
        2487 => x"13050900",
        2488 => x"ef000009",
        2489 => x"1305b400",
        2490 => x"93074400",
        2491 => x"137585ff",
        2492 => x"3307f540",
        2493 => x"e30cf5f8",
        2494 => x"3304e400",
        2495 => x"b387a740",
        2496 => x"2320f400",
        2497 => x"6ff09ff8",
        2498 => x"23a2e700",
        2499 => x"6ff05ffc",
        2500 => x"03274400",
        2501 => x"63968700",
        2502 => x"23a6e188",
        2503 => x"6ff01ffc",
        2504 => x"23a2e700",
        2505 => x"6ff09ffb",
        2506 => x"93070400",
        2507 => x"03244400",
        2508 => x"6ff09fec",
        2509 => x"13840700",
        2510 => x"83a74700",
        2511 => x"6ff01fee",
        2512 => x"93070700",
        2513 => x"6ff05ff2",
        2514 => x"9307c000",
        2515 => x"2320f900",
        2516 => x"13050900",
        2517 => x"ef00c001",
        2518 => x"6ff01ff3",
        2519 => x"23209500",
        2520 => x"6ff0dff7",
        2521 => x"23220000",
        2522 => x"73001000",
        2523 => x"67800000",
        2524 => x"67800000",
        2525 => x"130101fe",
        2526 => x"23282101",
        2527 => x"03a98500",
        2528 => x"232c8100",
        2529 => x"23263101",
        2530 => x"23225101",
        2531 => x"23206101",
        2532 => x"232e1100",
        2533 => x"232a9100",
        2534 => x"23244101",
        2535 => x"83aa0500",
        2536 => x"13840500",
        2537 => x"130b0600",
        2538 => x"93890600",
        2539 => x"63ec2609",
        2540 => x"8397c500",
        2541 => x"13f70748",
        2542 => x"63040708",
        2543 => x"03274401",
        2544 => x"93043000",
        2545 => x"83a50501",
        2546 => x"b384e402",
        2547 => x"13072000",
        2548 => x"b38aba40",
        2549 => x"130a0500",
        2550 => x"b3c4e402",
        2551 => x"13871600",
        2552 => x"33075701",
        2553 => x"63f4e400",
        2554 => x"93040700",
        2555 => x"93f70740",
        2556 => x"6386070a",
        2557 => x"93850400",
        2558 => x"13050a00",
        2559 => x"eff01fdb",
        2560 => x"13090500",
        2561 => x"630c050a",
        2562 => x"83250401",
        2563 => x"13860a00",
        2564 => x"efe05fb9",
        2565 => x"8357c400",
        2566 => x"93f7f7b7",
        2567 => x"93e70708",
        2568 => x"2316f400",
        2569 => x"23282401",
        2570 => x"232a9400",
        2571 => x"33095901",
        2572 => x"b3845441",
        2573 => x"23202401",
        2574 => x"23249400",
        2575 => x"13890900",
        2576 => x"63f42901",
        2577 => x"13890900",
        2578 => x"03250400",
        2579 => x"13060900",
        2580 => x"93050b00",
        2581 => x"efe05fb7",
        2582 => x"83278400",
        2583 => x"13050000",
        2584 => x"b3872741",
        2585 => x"2324f400",
        2586 => x"83270400",
        2587 => x"b3872701",
        2588 => x"2320f400",
        2589 => x"8320c101",
        2590 => x"03248101",
        2591 => x"83244101",
        2592 => x"03290101",
        2593 => x"8329c100",
        2594 => x"032a8100",
        2595 => x"832a4100",
        2596 => x"032b0100",
        2597 => x"13010102",
        2598 => x"67800000",
        2599 => x"13860400",
        2600 => x"13050a00",
        2601 => x"ef001060",
        2602 => x"13090500",
        2603 => x"e31c05f6",
        2604 => x"83250401",
        2605 => x"13050a00",
        2606 => x"eff09fb7",
        2607 => x"9307c000",
        2608 => x"2320fa00",
        2609 => x"8357c400",
        2610 => x"1305f0ff",
        2611 => x"93e70704",
        2612 => x"2316f400",
        2613 => x"6ff01ffa",
        2614 => x"83278600",
        2615 => x"130101fd",
        2616 => x"232e3101",
        2617 => x"23267101",
        2618 => x"23261102",
        2619 => x"23248102",
        2620 => x"23229102",
        2621 => x"23202103",
        2622 => x"232c4101",
        2623 => x"232a5101",
        2624 => x"23286101",
        2625 => x"23248101",
        2626 => x"23229101",
        2627 => x"2320a101",
        2628 => x"832b0600",
        2629 => x"93090600",
        2630 => x"63980712",
        2631 => x"13050000",
        2632 => x"8320c102",
        2633 => x"03248102",
        2634 => x"23a20900",
        2635 => x"83244102",
        2636 => x"03290102",
        2637 => x"8329c101",
        2638 => x"032a8101",
        2639 => x"832a4101",
        2640 => x"032b0101",
        2641 => x"832bc100",
        2642 => x"032c8100",
        2643 => x"832c4100",
        2644 => x"032d0100",
        2645 => x"13010103",
        2646 => x"67800000",
        2647 => x"03ab0b00",
        2648 => x"03ad4b00",
        2649 => x"938b8b00",
        2650 => x"03298400",
        2651 => x"832a0400",
        2652 => x"e3060dfe",
        2653 => x"63642d09",
        2654 => x"8317c400",
        2655 => x"13f70748",
        2656 => x"63020708",
        2657 => x"83244401",
        2658 => x"83250401",
        2659 => x"b3049c02",
        2660 => x"b38aba40",
        2661 => x"13871a00",
        2662 => x"3307a701",
        2663 => x"b3c49403",
        2664 => x"63f4e400",
        2665 => x"93040700",
        2666 => x"93f70740",
        2667 => x"638c070a",
        2668 => x"93850400",
        2669 => x"13050a00",
        2670 => x"eff05fbf",
        2671 => x"13090500",
        2672 => x"6302050c",
        2673 => x"83250401",
        2674 => x"13860a00",
        2675 => x"efe09f9d",
        2676 => x"8357c400",
        2677 => x"93f7f7b7",
        2678 => x"93e70708",
        2679 => x"2316f400",
        2680 => x"23282401",
        2681 => x"232a9400",
        2682 => x"33095901",
        2683 => x"b3845441",
        2684 => x"23202401",
        2685 => x"23249400",
        2686 => x"13090d00",
        2687 => x"63742d01",
        2688 => x"13090d00",
        2689 => x"03250400",
        2690 => x"93050b00",
        2691 => x"13060900",
        2692 => x"efe09f9b",
        2693 => x"83278400",
        2694 => x"330bab01",
        2695 => x"b3872741",
        2696 => x"2324f400",
        2697 => x"83270400",
        2698 => x"b3872701",
        2699 => x"2320f400",
        2700 => x"83a78900",
        2701 => x"b387a741",
        2702 => x"23a4f900",
        2703 => x"e38007ee",
        2704 => x"130d0000",
        2705 => x"6ff05ff2",
        2706 => x"130a0500",
        2707 => x"13840500",
        2708 => x"130b0000",
        2709 => x"130d0000",
        2710 => x"130c3000",
        2711 => x"930c2000",
        2712 => x"6ff09ff0",
        2713 => x"13860400",
        2714 => x"13050a00",
        2715 => x"ef009043",
        2716 => x"13090500",
        2717 => x"e31605f6",
        2718 => x"83250401",
        2719 => x"13050a00",
        2720 => x"eff01f9b",
        2721 => x"9307c000",
        2722 => x"2320fa00",
        2723 => x"8357c400",
        2724 => x"1305f0ff",
        2725 => x"93e70704",
        2726 => x"2316f400",
        2727 => x"23a40900",
        2728 => x"6ff01fe8",
        2729 => x"83d7c500",
        2730 => x"130101f5",
        2731 => x"2324810a",
        2732 => x"2322910a",
        2733 => x"2320210b",
        2734 => x"232c4109",
        2735 => x"2326110a",
        2736 => x"232e3109",
        2737 => x"232a5109",
        2738 => x"23286109",
        2739 => x"23267109",
        2740 => x"23248109",
        2741 => x"23229109",
        2742 => x"2320a109",
        2743 => x"232eb107",
        2744 => x"93f70708",
        2745 => x"130a0500",
        2746 => x"13890500",
        2747 => x"93040600",
        2748 => x"13840600",
        2749 => x"63880706",
        2750 => x"83a70501",
        2751 => x"63940706",
        2752 => x"93050004",
        2753 => x"eff09faa",
        2754 => x"2320a900",
        2755 => x"2328a900",
        2756 => x"63160504",
        2757 => x"9307c000",
        2758 => x"2320fa00",
        2759 => x"1305f0ff",
        2760 => x"8320c10a",
        2761 => x"0324810a",
        2762 => x"8324410a",
        2763 => x"0329010a",
        2764 => x"8329c109",
        2765 => x"032a8109",
        2766 => x"832a4109",
        2767 => x"032b0109",
        2768 => x"832bc108",
        2769 => x"032c8108",
        2770 => x"832c4108",
        2771 => x"032d0108",
        2772 => x"832dc107",
        2773 => x"1301010b",
        2774 => x"67800000",
        2775 => x"93070004",
        2776 => x"232af900",
        2777 => x"93070002",
        2778 => x"a304f102",
        2779 => x"93070003",
        2780 => x"23220102",
        2781 => x"2305f102",
        2782 => x"23268100",
        2783 => x"930c5002",
        2784 => x"374b0000",
        2785 => x"b74b0000",
        2786 => x"374d0000",
        2787 => x"372c0000",
        2788 => x"930a0000",
        2789 => x"13840400",
        2790 => x"83470400",
        2791 => x"63840700",
        2792 => x"639c970d",
        2793 => x"b30d9440",
        2794 => x"63069402",
        2795 => x"93860d00",
        2796 => x"13860400",
        2797 => x"93050900",
        2798 => x"13050a00",
        2799 => x"eff09fbb",
        2800 => x"9307f0ff",
        2801 => x"6304f524",
        2802 => x"83274102",
        2803 => x"b387b701",
        2804 => x"2322f102",
        2805 => x"83470400",
        2806 => x"638a0722",
        2807 => x"9307f0ff",
        2808 => x"93041400",
        2809 => x"23280100",
        2810 => x"232e0100",
        2811 => x"232af100",
        2812 => x"232c0100",
        2813 => x"a3090104",
        2814 => x"23240106",
        2815 => x"930d1000",
        2816 => x"83c50400",
        2817 => x"13065000",
        2818 => x"1305cbba",
        2819 => x"ef00101e",
        2820 => x"83270101",
        2821 => x"13841400",
        2822 => x"63140506",
        2823 => x"13f70701",
        2824 => x"63060700",
        2825 => x"13070002",
        2826 => x"a309e104",
        2827 => x"13f78700",
        2828 => x"63060700",
        2829 => x"1307b002",
        2830 => x"a309e104",
        2831 => x"83c60400",
        2832 => x"1307a002",
        2833 => x"638ce604",
        2834 => x"8327c101",
        2835 => x"13840400",
        2836 => x"93060000",
        2837 => x"13069000",
        2838 => x"1305a000",
        2839 => x"03470400",
        2840 => x"93051400",
        2841 => x"130707fd",
        2842 => x"637ee608",
        2843 => x"63840604",
        2844 => x"232ef100",
        2845 => x"6f000004",
        2846 => x"13041400",
        2847 => x"6ff0dff1",
        2848 => x"1307cbba",
        2849 => x"3305e540",
        2850 => x"3395ad00",
        2851 => x"b3e7a700",
        2852 => x"2328f100",
        2853 => x"93040400",
        2854 => x"6ff09ff6",
        2855 => x"0327c100",
        2856 => x"93064700",
        2857 => x"03270700",
        2858 => x"2326d100",
        2859 => x"63420704",
        2860 => x"232ee100",
        2861 => x"03470400",
        2862 => x"9307e002",
        2863 => x"6314f708",
        2864 => x"03471400",
        2865 => x"9307a002",
        2866 => x"6318f704",
        2867 => x"8327c100",
        2868 => x"13042400",
        2869 => x"13874700",
        2870 => x"83a70700",
        2871 => x"2326e100",
        2872 => x"63d40700",
        2873 => x"9307f0ff",
        2874 => x"232af100",
        2875 => x"6f008005",
        2876 => x"3307e040",
        2877 => x"93e72700",
        2878 => x"232ee100",
        2879 => x"2328f100",
        2880 => x"6ff05ffb",
        2881 => x"b387a702",
        2882 => x"13840500",
        2883 => x"93061000",
        2884 => x"b387e700",
        2885 => x"6ff09ff4",
        2886 => x"13041400",
        2887 => x"232a0100",
        2888 => x"93060000",
        2889 => x"93070000",
        2890 => x"13069000",
        2891 => x"1305a000",
        2892 => x"03470400",
        2893 => x"93051400",
        2894 => x"130707fd",
        2895 => x"6372e608",
        2896 => x"e39406fa",
        2897 => x"83450400",
        2898 => x"13063000",
        2899 => x"13854bbb",
        2900 => x"ef00d009",
        2901 => x"63020502",
        2902 => x"93874bbb",
        2903 => x"3305f540",
        2904 => x"83270101",
        2905 => x"13070004",
        2906 => x"3317a700",
        2907 => x"b3e7e700",
        2908 => x"13041400",
        2909 => x"2328f100",
        2910 => x"83450400",
        2911 => x"13066000",
        2912 => x"13058dbb",
        2913 => x"93041400",
        2914 => x"2304b102",
        2915 => x"ef001006",
        2916 => x"63080508",
        2917 => x"63980a04",
        2918 => x"03270101",
        2919 => x"8327c100",
        2920 => x"13770710",
        2921 => x"63080702",
        2922 => x"93874700",
        2923 => x"2326f100",
        2924 => x"83274102",
        2925 => x"b3873701",
        2926 => x"2322f102",
        2927 => x"6ff09fdd",
        2928 => x"b387a702",
        2929 => x"13840500",
        2930 => x"93061000",
        2931 => x"b387e700",
        2932 => x"6ff01ff6",
        2933 => x"93877700",
        2934 => x"93f787ff",
        2935 => x"93878700",
        2936 => x"6ff0dffc",
        2937 => x"1307c100",
        2938 => x"93064c77",
        2939 => x"13060900",
        2940 => x"93050101",
        2941 => x"13050a00",
        2942 => x"97000000",
        2943 => x"e7000000",
        2944 => x"9307f0ff",
        2945 => x"93090500",
        2946 => x"e314f5fa",
        2947 => x"8357c900",
        2948 => x"93f70704",
        2949 => x"e39407d0",
        2950 => x"03254102",
        2951 => x"6ff05fd0",
        2952 => x"1307c100",
        2953 => x"93064c77",
        2954 => x"13060900",
        2955 => x"93050101",
        2956 => x"13050a00",
        2957 => x"ef00801b",
        2958 => x"6ff09ffc",
        2959 => x"130101fd",
        2960 => x"232a5101",
        2961 => x"83a70501",
        2962 => x"930a0700",
        2963 => x"03a78500",
        2964 => x"23248102",
        2965 => x"23202103",
        2966 => x"232e3101",
        2967 => x"232c4101",
        2968 => x"23261102",
        2969 => x"23229102",
        2970 => x"23286101",
        2971 => x"23267101",
        2972 => x"93090500",
        2973 => x"13840500",
        2974 => x"13090600",
        2975 => x"138a0600",
        2976 => x"63d4e700",
        2977 => x"93070700",
        2978 => x"2320f900",
        2979 => x"03473404",
        2980 => x"63060700",
        2981 => x"93871700",
        2982 => x"2320f900",
        2983 => x"83270400",
        2984 => x"93f70702",
        2985 => x"63880700",
        2986 => x"83270900",
        2987 => x"93872700",
        2988 => x"2320f900",
        2989 => x"83240400",
        2990 => x"93f46400",
        2991 => x"639e0400",
        2992 => x"130b9401",
        2993 => x"930bf0ff",
        2994 => x"8327c400",
        2995 => x"03270900",
        2996 => x"b387e740",
        2997 => x"63c2f408",
        2998 => x"83473404",
        2999 => x"b336f000",
        3000 => x"83270400",
        3001 => x"93f70702",
        3002 => x"6390070c",
        3003 => x"13063404",
        3004 => x"93050a00",
        3005 => x"13850900",
        3006 => x"e7800a00",
        3007 => x"9307f0ff",
        3008 => x"6308f506",
        3009 => x"83270400",
        3010 => x"13074000",
        3011 => x"93040000",
        3012 => x"93f76700",
        3013 => x"639ce700",
        3014 => x"8324c400",
        3015 => x"83270900",
        3016 => x"b384f440",
        3017 => x"63d40400",
        3018 => x"93040000",
        3019 => x"83278400",
        3020 => x"03270401",
        3021 => x"6356f700",
        3022 => x"b387e740",
        3023 => x"b384f400",
        3024 => x"13090000",
        3025 => x"1304a401",
        3026 => x"130bf0ff",
        3027 => x"63902409",
        3028 => x"13050000",
        3029 => x"6f000002",
        3030 => x"93061000",
        3031 => x"13060b00",
        3032 => x"93050a00",
        3033 => x"13850900",
        3034 => x"e7800a00",
        3035 => x"631a7503",
        3036 => x"1305f0ff",
        3037 => x"8320c102",
        3038 => x"03248102",
        3039 => x"83244102",
        3040 => x"03290102",
        3041 => x"8329c101",
        3042 => x"032a8101",
        3043 => x"832a4101",
        3044 => x"032b0101",
        3045 => x"832bc100",
        3046 => x"13010103",
        3047 => x"67800000",
        3048 => x"93841400",
        3049 => x"6ff05ff2",
        3050 => x"3307d400",
        3051 => x"13060003",
        3052 => x"a301c704",
        3053 => x"03475404",
        3054 => x"93871600",
        3055 => x"b307f400",
        3056 => x"93862600",
        3057 => x"a381e704",
        3058 => x"6ff05ff2",
        3059 => x"93061000",
        3060 => x"13060400",
        3061 => x"93050a00",
        3062 => x"13850900",
        3063 => x"e7800a00",
        3064 => x"e30865f9",
        3065 => x"13091900",
        3066 => x"6ff05ff6",
        3067 => x"130101fd",
        3068 => x"23248102",
        3069 => x"23202103",
        3070 => x"232e3101",
        3071 => x"232c4101",
        3072 => x"23261102",
        3073 => x"23229102",
        3074 => x"232a5101",
        3075 => x"23286101",
        3076 => x"138a0600",
        3077 => x"83c68501",
        3078 => x"93078007",
        3079 => x"13090500",
        3080 => x"13840500",
        3081 => x"93090600",
        3082 => x"63eed700",
        3083 => x"93072006",
        3084 => x"13863504",
        3085 => x"63eed700",
        3086 => x"63840628",
        3087 => x"93078005",
        3088 => x"6380f622",
        3089 => x"93042404",
        3090 => x"2301d404",
        3091 => x"6f004004",
        3092 => x"9387d6f9",
        3093 => x"93f7f70f",
        3094 => x"93055001",
        3095 => x"e3e4f5fe",
        3096 => x"b7450000",
        3097 => x"93972700",
        3098 => x"938585be",
        3099 => x"b387b700",
        3100 => x"83a70700",
        3101 => x"67800700",
        3102 => x"83270700",
        3103 => x"93042404",
        3104 => x"93864700",
        3105 => x"83a70700",
        3106 => x"2320d700",
        3107 => x"2301f404",
        3108 => x"93071000",
        3109 => x"6f008026",
        3110 => x"83270400",
        3111 => x"03250700",
        3112 => x"93f60708",
        3113 => x"93054500",
        3114 => x"63860602",
        3115 => x"83270500",
        3116 => x"2320b700",
        3117 => x"37480000",
        3118 => x"63d80700",
        3119 => x"1307d002",
        3120 => x"b307f040",
        3121 => x"a301e404",
        3122 => x"130808bc",
        3123 => x"1307a000",
        3124 => x"6f004006",
        3125 => x"93f60704",
        3126 => x"83270500",
        3127 => x"2320b700",
        3128 => x"e38a06fc",
        3129 => x"93970701",
        3130 => x"93d70741",
        3131 => x"6ff09ffc",
        3132 => x"03250400",
        3133 => x"83250700",
        3134 => x"13780508",
        3135 => x"83a70500",
        3136 => x"93854500",
        3137 => x"631a0800",
        3138 => x"13750504",
        3139 => x"63060500",
        3140 => x"93970701",
        3141 => x"93d70701",
        3142 => x"2320b700",
        3143 => x"37480000",
        3144 => x"1307f006",
        3145 => x"130808bc",
        3146 => x"639ae614",
        3147 => x"13078000",
        3148 => x"a3010404",
        3149 => x"83264400",
        3150 => x"2324d400",
        3151 => x"63ce0600",
        3152 => x"83250400",
        3153 => x"b3e6d700",
        3154 => x"93040600",
        3155 => x"93f5b5ff",
        3156 => x"2320b400",
        3157 => x"63840602",
        3158 => x"93040600",
        3159 => x"b3f6e702",
        3160 => x"9384f4ff",
        3161 => x"b306d800",
        3162 => x"83c60600",
        3163 => x"2380d400",
        3164 => x"93860700",
        3165 => x"b3d7e702",
        3166 => x"e3f2e6fe",
        3167 => x"93078000",
        3168 => x"6314f702",
        3169 => x"83270400",
        3170 => x"93f71700",
        3171 => x"638e0700",
        3172 => x"03274400",
        3173 => x"83270401",
        3174 => x"63c8e700",
        3175 => x"93070003",
        3176 => x"a38ff4fe",
        3177 => x"9384f4ff",
        3178 => x"33069640",
        3179 => x"2328c400",
        3180 => x"13070a00",
        3181 => x"93860900",
        3182 => x"1306c100",
        3183 => x"93050400",
        3184 => x"13050900",
        3185 => x"eff09fc7",
        3186 => x"930af0ff",
        3187 => x"631e5513",
        3188 => x"1305f0ff",
        3189 => x"8320c102",
        3190 => x"03248102",
        3191 => x"83244102",
        3192 => x"03290102",
        3193 => x"8329c101",
        3194 => x"032a8101",
        3195 => x"832a4101",
        3196 => x"032b0101",
        3197 => x"13010103",
        3198 => x"67800000",
        3199 => x"83270400",
        3200 => x"93e70702",
        3201 => x"2320f400",
        3202 => x"37480000",
        3203 => x"93068007",
        3204 => x"130848bd",
        3205 => x"a302d404",
        3206 => x"83260400",
        3207 => x"83250700",
        3208 => x"13f50608",
        3209 => x"83a70500",
        3210 => x"93854500",
        3211 => x"631a0500",
        3212 => x"13f50604",
        3213 => x"63060500",
        3214 => x"93970701",
        3215 => x"93d70701",
        3216 => x"2320b700",
        3217 => x"13f71600",
        3218 => x"63060700",
        3219 => x"93e60602",
        3220 => x"2320d400",
        3221 => x"638c0700",
        3222 => x"13070001",
        3223 => x"6ff05fed",
        3224 => x"37480000",
        3225 => x"130808bc",
        3226 => x"6ff0dffa",
        3227 => x"03270400",
        3228 => x"1377f7fd",
        3229 => x"2320e400",
        3230 => x"6ff01ffe",
        3231 => x"1307a000",
        3232 => x"6ff01feb",
        3233 => x"83260400",
        3234 => x"83270700",
        3235 => x"83254401",
        3236 => x"13f80608",
        3237 => x"13854700",
        3238 => x"630a0800",
        3239 => x"2320a700",
        3240 => x"83a70700",
        3241 => x"23a0b700",
        3242 => x"6f008001",
        3243 => x"2320a700",
        3244 => x"93f60604",
        3245 => x"83a70700",
        3246 => x"e38606fe",
        3247 => x"2390b700",
        3248 => x"23280400",
        3249 => x"93040600",
        3250 => x"6ff09fee",
        3251 => x"83270700",
        3252 => x"03264400",
        3253 => x"93050000",
        3254 => x"93864700",
        3255 => x"2320d700",
        3256 => x"83a40700",
        3257 => x"13850400",
        3258 => x"ef004030",
        3259 => x"63060500",
        3260 => x"33059540",
        3261 => x"2322a400",
        3262 => x"83274400",
        3263 => x"2328f400",
        3264 => x"a3010404",
        3265 => x"6ff0dfea",
        3266 => x"83260401",
        3267 => x"13860400",
        3268 => x"93850900",
        3269 => x"13050900",
        3270 => x"e7000a00",
        3271 => x"e30a55eb",
        3272 => x"83270400",
        3273 => x"93f72700",
        3274 => x"63940704",
        3275 => x"8327c100",
        3276 => x"0325c400",
        3277 => x"e350f5ea",
        3278 => x"13850700",
        3279 => x"6ff09fe9",
        3280 => x"93061000",
        3281 => x"13860a00",
        3282 => x"93850900",
        3283 => x"13050900",
        3284 => x"e7000a00",
        3285 => x"e30e65e7",
        3286 => x"93841400",
        3287 => x"8327c400",
        3288 => x"0327c100",
        3289 => x"b387e740",
        3290 => x"e3ccf4fc",
        3291 => x"6ff01ffc",
        3292 => x"93040000",
        3293 => x"930a9401",
        3294 => x"130bf0ff",
        3295 => x"6ff01ffe",
        3296 => x"8397c500",
        3297 => x"130101fe",
        3298 => x"232c8100",
        3299 => x"232a9100",
        3300 => x"232e1100",
        3301 => x"23282101",
        3302 => x"23263101",
        3303 => x"13f78700",
        3304 => x"93040500",
        3305 => x"13840500",
        3306 => x"631a0712",
        3307 => x"03a74500",
        3308 => x"6346e000",
        3309 => x"03a70504",
        3310 => x"6356e010",
        3311 => x"0327c402",
        3312 => x"63020710",
        3313 => x"03a90400",
        3314 => x"93963701",
        3315 => x"23a00400",
        3316 => x"83250402",
        3317 => x"63dc060a",
        3318 => x"03264405",
        3319 => x"8357c400",
        3320 => x"93f74700",
        3321 => x"638e0700",
        3322 => x"83274400",
        3323 => x"3306f640",
        3324 => x"83274403",
        3325 => x"63860700",
        3326 => x"83270404",
        3327 => x"3306f640",
        3328 => x"8327c402",
        3329 => x"83250402",
        3330 => x"93060000",
        3331 => x"13850400",
        3332 => x"e7800700",
        3333 => x"1307f0ff",
        3334 => x"8357c400",
        3335 => x"6312e502",
        3336 => x"83a60400",
        3337 => x"1307d001",
        3338 => x"6362d70a",
        3339 => x"37074020",
        3340 => x"13071700",
        3341 => x"3357d700",
        3342 => x"13771700",
        3343 => x"63080708",
        3344 => x"03270401",
        3345 => x"23220400",
        3346 => x"2320e400",
        3347 => x"13973701",
        3348 => x"635c0700",
        3349 => x"9307f0ff",
        3350 => x"6316f500",
        3351 => x"83a70400",
        3352 => x"63940700",
        3353 => x"232aa404",
        3354 => x"83254403",
        3355 => x"23a02401",
        3356 => x"638a0504",
        3357 => x"93074404",
        3358 => x"6386f500",
        3359 => x"13850400",
        3360 => x"efe01ffb",
        3361 => x"232a0402",
        3362 => x"6f00c003",
        3363 => x"13060000",
        3364 => x"93061000",
        3365 => x"13850400",
        3366 => x"e7000700",
        3367 => x"9307f0ff",
        3368 => x"13060500",
        3369 => x"e31cf5f2",
        3370 => x"83a70400",
        3371 => x"e38807f2",
        3372 => x"1307d001",
        3373 => x"6386e700",
        3374 => x"13076001",
        3375 => x"6394e706",
        3376 => x"23a02401",
        3377 => x"13050000",
        3378 => x"6f00c006",
        3379 => x"93e70704",
        3380 => x"93970701",
        3381 => x"93d70741",
        3382 => x"6f004005",
        3383 => x"83a90501",
        3384 => x"e38209fe",
        3385 => x"03a90500",
        3386 => x"93f73700",
        3387 => x"23a03501",
        3388 => x"33093941",
        3389 => x"13070000",
        3390 => x"63940700",
        3391 => x"03a74501",
        3392 => x"2324e400",
        3393 => x"e35020fd",
        3394 => x"83278402",
        3395 => x"83250402",
        3396 => x"93060900",
        3397 => x"13860900",
        3398 => x"13850400",
        3399 => x"e7800700",
        3400 => x"6348a002",
        3401 => x"8317c400",
        3402 => x"93e70704",
        3403 => x"2316f400",
        3404 => x"1305f0ff",
        3405 => x"8320c101",
        3406 => x"03248101",
        3407 => x"83244101",
        3408 => x"03290101",
        3409 => x"8329c100",
        3410 => x"13010102",
        3411 => x"67800000",
        3412 => x"b389a900",
        3413 => x"3309a940",
        3414 => x"6ff0dffa",
        3415 => x"83a70501",
        3416 => x"638e0704",
        3417 => x"130101fe",
        3418 => x"232c8100",
        3419 => x"232e1100",
        3420 => x"13040500",
        3421 => x"630c0500",
        3422 => x"83270502",
        3423 => x"63980700",
        3424 => x"2326b100",
        3425 => x"efe05f85",
        3426 => x"8325c100",
        3427 => x"8397c500",
        3428 => x"638c0700",
        3429 => x"13050400",
        3430 => x"03248101",
        3431 => x"8320c101",
        3432 => x"13010102",
        3433 => x"6ff0dfdd",
        3434 => x"8320c101",
        3435 => x"03248101",
        3436 => x"13050000",
        3437 => x"13010102",
        3438 => x"67800000",
        3439 => x"13050000",
        3440 => x"67800000",
        3441 => x"93050500",
        3442 => x"631e0500",
        3443 => x"b7350000",
        3444 => x"37050020",
        3445 => x"13868181",
        3446 => x"9385c555",
        3447 => x"13054502",
        3448 => x"6fe0df84",
        3449 => x"03a54187",
        3450 => x"6ff05ff7",
        3451 => x"93f5f50f",
        3452 => x"3306c500",
        3453 => x"6316c500",
        3454 => x"13050000",
        3455 => x"67800000",
        3456 => x"83470500",
        3457 => x"e38cb7fe",
        3458 => x"13051500",
        3459 => x"6ff09ffe",
        3460 => x"130101ff",
        3461 => x"23248100",
        3462 => x"23229100",
        3463 => x"13040500",
        3464 => x"13850500",
        3465 => x"93050600",
        3466 => x"23261100",
        3467 => x"23a20188",
        3468 => x"efd09fdd",
        3469 => x"9307f0ff",
        3470 => x"6318f500",
        3471 => x"83a74188",
        3472 => x"63840700",
        3473 => x"2320f400",
        3474 => x"8320c100",
        3475 => x"03248100",
        3476 => x"83244100",
        3477 => x"13010101",
        3478 => x"67800000",
        3479 => x"130101ff",
        3480 => x"23248100",
        3481 => x"23229100",
        3482 => x"13040500",
        3483 => x"13850500",
        3484 => x"23261100",
        3485 => x"23a20188",
        3486 => x"efe0cf80",
        3487 => x"9307f0ff",
        3488 => x"6318f500",
        3489 => x"83a74188",
        3490 => x"63840700",
        3491 => x"2320f400",
        3492 => x"8320c100",
        3493 => x"03248100",
        3494 => x"83244100",
        3495 => x"13010101",
        3496 => x"67800000",
        3497 => x"130101fe",
        3498 => x"232c8100",
        3499 => x"232e1100",
        3500 => x"232a9100",
        3501 => x"23282101",
        3502 => x"23263101",
        3503 => x"23244101",
        3504 => x"13040600",
        3505 => x"63940502",
        3506 => x"03248101",
        3507 => x"8320c101",
        3508 => x"83244101",
        3509 => x"03290101",
        3510 => x"8329c100",
        3511 => x"032a8100",
        3512 => x"93050600",
        3513 => x"13010102",
        3514 => x"6fe05fec",
        3515 => x"63180602",
        3516 => x"efe01fd4",
        3517 => x"93040000",
        3518 => x"8320c101",
        3519 => x"03248101",
        3520 => x"03290101",
        3521 => x"8329c100",
        3522 => x"032a8100",
        3523 => x"13850400",
        3524 => x"83244101",
        3525 => x"13010102",
        3526 => x"67800000",
        3527 => x"130a0500",
        3528 => x"93840500",
        3529 => x"ef008005",
        3530 => x"13090500",
        3531 => x"63668500",
        3532 => x"93571500",
        3533 => x"e3e287fc",
        3534 => x"93050400",
        3535 => x"13050a00",
        3536 => x"efe0dfe6",
        3537 => x"93090500",
        3538 => x"63160500",
        3539 => x"93840900",
        3540 => x"6ff09ffa",
        3541 => x"13060400",
        3542 => x"63748900",
        3543 => x"13060900",
        3544 => x"93850400",
        3545 => x"13850900",
        3546 => x"efd0dfc3",
        3547 => x"93850400",
        3548 => x"13050a00",
        3549 => x"efe0dfcb",
        3550 => x"6ff05ffd",
        3551 => x"83a7c5ff",
        3552 => x"1385c7ff",
        3553 => x"63d80700",
        3554 => x"b385a500",
        3555 => x"83a70500",
        3556 => x"3305f500",
        3557 => x"67800000",
        3558 => x"10000000",
        3559 => x"00000000",
        3560 => x"037a5200",
        3561 => x"017c0101",
        3562 => x"1b0d0200",
        3563 => x"10000000",
        3564 => x"18000000",
        3565 => x"48cfffff",
        3566 => x"78040000",
        3567 => x"00000000",
        3568 => x"10000000",
        3569 => x"00000000",
        3570 => x"037a5200",
        3571 => x"017c0101",
        3572 => x"1b0d0200",
        3573 => x"10000000",
        3574 => x"18000000",
        3575 => x"98d3ffff",
        3576 => x"30040000",
        3577 => x"00000000",
        3578 => x"10000000",
        3579 => x"00000000",
        3580 => x"037a5200",
        3581 => x"017c0101",
        3582 => x"1b0d0200",
        3583 => x"10000000",
        3584 => x"18000000",
        3585 => x"a0d7ffff",
        3586 => x"e4030000",
        3587 => x"00000000",
        3588 => x"30313233",
        3589 => x"34353637",
        3590 => x"38396162",
        3591 => x"63646566",
        3592 => x"00000000",
        3593 => x"a4040000",
        3594 => x"dc030000",
        3595 => x"dc030000",
        3596 => x"dc030000",
        3597 => x"b0040000",
        3598 => x"dc030000",
        3599 => x"dc030000",
        3600 => x"dc030000",
        3601 => x"dc030000",
        3602 => x"dc030000",
        3603 => x"dc030000",
        3604 => x"dc030000",
        3605 => x"dc030000",
        3606 => x"dc030000",
        3607 => x"dc030000",
        3608 => x"bc040000",
        3609 => x"dc030000",
        3610 => x"c8040000",
        3611 => x"d4040000",
        3612 => x"dc030000",
        3613 => x"e0040000",
        3614 => x"ec040000",
        3615 => x"dc030000",
        3616 => x"f8040000",
        3617 => x"98040000",
        3618 => x"dc030000",
        3619 => x"dc030000",
        3620 => x"dc030000",
        3621 => x"04050000",
        3622 => x"dc030000",
        3623 => x"dc030000",
        3624 => x"dc030000",
        3625 => x"dc030000",
        3626 => x"dc030000",
        3627 => x"dc030000",
        3628 => x"dc030000",
        3629 => x"14050000",
        3630 => x"a8050000",
        3631 => x"c0050000",
        3632 => x"f0050000",
        3633 => x"70050000",
        3634 => x"70050000",
        3635 => x"70050000",
        3636 => x"70050000",
        3637 => x"70050000",
        3638 => x"70050000",
        3639 => x"d8050000",
        3640 => x"70050000",
        3641 => x"70050000",
        3642 => x"70050000",
        3643 => x"70050000",
        3644 => x"88050000",
        3645 => x"88050000",
        3646 => x"a8050000",
        3647 => x"70050000",
        3648 => x"70050000",
        3649 => x"70050000",
        3650 => x"70050000",
        3651 => x"9c050000",
        3652 => x"08060000",
        3653 => x"30060000",
        3654 => x"70050000",
        3655 => x"70050000",
        3656 => x"70050000",
        3657 => x"70050000",
        3658 => x"70050000",
        3659 => x"70050000",
        3660 => x"70050000",
        3661 => x"70050000",
        3662 => x"70050000",
        3663 => x"70050000",
        3664 => x"70050000",
        3665 => x"70050000",
        3666 => x"70050000",
        3667 => x"70050000",
        3668 => x"88050000",
        3669 => x"88050000",
        3670 => x"70050000",
        3671 => x"70050000",
        3672 => x"70050000",
        3673 => x"70050000",
        3674 => x"70050000",
        3675 => x"70050000",
        3676 => x"70050000",
        3677 => x"70050000",
        3678 => x"70050000",
        3679 => x"70050000",
        3680 => x"70050000",
        3681 => x"70050000",
        3682 => x"9c050000",
        3683 => x"00010202",
        3684 => x"03030303",
        3685 => x"04040404",
        3686 => x"04040404",
        3687 => x"05050505",
        3688 => x"05050505",
        3689 => x"05050505",
        3690 => x"05050505",
        3691 => x"06060606",
        3692 => x"06060606",
        3693 => x"06060606",
        3694 => x"06060606",
        3695 => x"06060606",
        3696 => x"06060606",
        3697 => x"06060606",
        3698 => x"06060606",
        3699 => x"07070707",
        3700 => x"07070707",
        3701 => x"07070707",
        3702 => x"07070707",
        3703 => x"07070707",
        3704 => x"07070707",
        3705 => x"07070707",
        3706 => x"07070707",
        3707 => x"07070707",
        3708 => x"07070707",
        3709 => x"07070707",
        3710 => x"07070707",
        3711 => x"07070707",
        3712 => x"07070707",
        3713 => x"07070707",
        3714 => x"07070707",
        3715 => x"08080808",
        3716 => x"08080808",
        3717 => x"08080808",
        3718 => x"08080808",
        3719 => x"08080808",
        3720 => x"08080808",
        3721 => x"08080808",
        3722 => x"08080808",
        3723 => x"08080808",
        3724 => x"08080808",
        3725 => x"08080808",
        3726 => x"08080808",
        3727 => x"08080808",
        3728 => x"08080808",
        3729 => x"08080808",
        3730 => x"08080808",
        3731 => x"08080808",
        3732 => x"08080808",
        3733 => x"08080808",
        3734 => x"08080808",
        3735 => x"08080808",
        3736 => x"08080808",
        3737 => x"08080808",
        3738 => x"08080808",
        3739 => x"08080808",
        3740 => x"08080808",
        3741 => x"08080808",
        3742 => x"08080808",
        3743 => x"08080808",
        3744 => x"08080808",
        3745 => x"08080808",
        3746 => x"08080808",
        3747 => x"0d0a4542",
        3748 => x"5245414b",
        3749 => x"21206d65",
        3750 => x"7063203d",
        3751 => x"20000000",
        3752 => x"20696e73",
        3753 => x"6e203d20",
        3754 => x"00000000",
        3755 => x"0d0a0000",
        3756 => x"0d0a0a44",
        3757 => x"6973706c",
        3758 => x"6179696e",
        3759 => x"67207468",
        3760 => x"65207469",
        3761 => x"6d652070",
        3762 => x"61737365",
        3763 => x"64207369",
        3764 => x"6e636520",
        3765 => x"72657365",
        3766 => x"740d0a0a",
        3767 => x"00000000",
        3768 => x"2530356c",
        3769 => x"643a2530",
        3770 => x"366c6420",
        3771 => x"20202530",
        3772 => x"326c643a",
        3773 => x"2530326c",
        3774 => x"643a2530",
        3775 => x"326c640d",
        3776 => x"00000000",
        3777 => x"696e7465",
        3778 => x"72727570",
        3779 => x"745f6469",
        3780 => x"72656374",
        3781 => x"00000000",
        3782 => x"54485541",
        3783 => x"53205249",
        3784 => x"53432d56",
        3785 => x"20525633",
        3786 => x"32494d20",
        3787 => x"62617265",
        3788 => x"206d6574",
        3789 => x"616c2070",
        3790 => x"726f6365",
        3791 => x"73736f72",
        3792 => x"00000000",
        3793 => x"54686520",
        3794 => x"48616775",
        3795 => x"6520556e",
        3796 => x"69766572",
        3797 => x"73697479",
        3798 => x"206f6620",
        3799 => x"4170706c",
        3800 => x"69656420",
        3801 => x"53636965",
        3802 => x"6e636573",
        3803 => x"00000000",
        3804 => x"44657061",
        3805 => x"72746d65",
        3806 => x"6e74206f",
        3807 => x"6620456c",
        3808 => x"65637472",
        3809 => x"6963616c",
        3810 => x"20456e67",
        3811 => x"696e6565",
        3812 => x"72696e67",
        3813 => x"00000000",
        3814 => x"4a2e452e",
        3815 => x"4a2e206f",
        3816 => x"70206465",
        3817 => x"6e204272",
        3818 => x"6f757700",
        3819 => x"232d302b",
        3820 => x"20000000",
        3821 => x"686c4c00",
        3822 => x"65666745",
        3823 => x"46470000",
        3824 => x"30313233",
        3825 => x"34353637",
        3826 => x"38394142",
        3827 => x"43444546",
        3828 => x"00000000",
        3829 => x"30313233",
        3830 => x"34353637",
        3831 => x"38396162",
        3832 => x"63646566",
        3833 => x"00000000",
        3834 => x"78300000",
        3835 => x"98300000",
        3836 => x"44300000",
        3837 => x"44300000",
        3838 => x"44300000",
        3839 => x"44300000",
        3840 => x"98300000",
        3841 => x"44300000",
        3842 => x"44300000",
        3843 => x"44300000",
        3844 => x"44300000",
        3845 => x"84320000",
        3846 => x"f0300000",
        3847 => x"fc310000",
        3848 => x"44300000",
        3849 => x"44300000",
        3850 => x"cc320000",
        3851 => x"44300000",
        3852 => x"f0300000",
        3853 => x"44300000",
        3854 => x"44300000",
        3855 => x"08320000",
        3856 => x"043b0000",
        3857 => x"183b0000",
        3858 => x"443b0000",
        3859 => x"703b0000",
        3860 => x"983b0000",
        3861 => x"00000000",
        3862 => x"00000000",
        3863 => x"03000000",
        3864 => x"90000020",
        3865 => x"00000000",
        3866 => x"90000020",
        3867 => x"f8000020",
        3868 => x"60010020",
        3869 => x"00000000",
        3870 => x"00000000",
        3871 => x"00000000",
        3872 => x"00000000",
        3873 => x"00000000",
        3874 => x"00000000",
        3875 => x"00000000",
        3876 => x"00000000",
        3877 => x"00000000",
        3878 => x"00000000",
        3879 => x"00000000",
        3880 => x"00000000",
        3881 => x"00000000",
        3882 => x"00000000",
        3883 => x"00000000",
        3884 => x"78000020",
        3885 => x"24000020",
        3886 => x"00000000"
            );
end package rom_image;
