-- srec2vhdl table generator
-- for input file 'bootloader.srec'
-- date: Mon Apr 29 18:20:12 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package bootrom_image is
    constant bootrom_contents : memory_type := (
           0 => x"97020000",
           1 => x"93828264",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"b7070020",
           9 => x"93870700",
          10 => x"13070500",
          11 => x"3386e740",
          12 => x"63f4e700",
          13 => x"13060000",
          14 => x"93050000",
          15 => x"13050500",
          16 => x"ef00c060",
          17 => x"37050020",
          18 => x"b7070020",
          19 => x"93870700",
          20 => x"13070500",
          21 => x"3386e740",
          22 => x"63f4e700",
          23 => x"13060000",
          24 => x"b7150010",
          25 => x"9385c5f1",
          26 => x"13050500",
          27 => x"ef00c05f",
          28 => x"ef001030",
          29 => x"37c50100",
          30 => x"93051000",
          31 => x"13050520",
          32 => x"ef00c07e",
          33 => x"37150010",
          34 => x"130585db",
          35 => x"ef00d002",
          36 => x"37150010",
          37 => x"1305c5dd",
          38 => x"ef001002",
          39 => x"732510fc",
          40 => x"37190010",
          41 => x"ef00101d",
          42 => x"130589dd",
          43 => x"ef00d000",
          44 => x"b70700f0",
          45 => x"1307f03f",
          46 => x"370a1000",
          47 => x"b709a000",
          48 => x"23a2e700",
          49 => x"93041000",
          50 => x"130afaff",
          51 => x"b70a00f0",
          52 => x"93891900",
          53 => x"b3f74401",
          54 => x"639c0700",
          55 => x"1305a002",
          56 => x"ef00807b",
          57 => x"83a74a00",
          58 => x"93d71700",
          59 => x"23a2fa00",
          60 => x"ef00c05b",
          61 => x"13040500",
          62 => x"63160504",
          63 => x"93841400",
          64 => x"e39a34fd",
          65 => x"b70700f0",
          66 => x"23a20700",
          67 => x"631a0400",
          68 => x"93050000",
          69 => x"13050000",
          70 => x"ef004075",
          71 => x"e7000400",
          72 => x"ef00c059",
          73 => x"1375f50f",
          74 => x"93071002",
          75 => x"6300f502",
          76 => x"93074002",
          77 => x"93040000",
          78 => x"6316f520",
          79 => x"13041000",
          80 => x"6f00c001",
          81 => x"13041000",
          82 => x"6ff0dffb",
          83 => x"37150010",
          84 => x"130505df",
          85 => x"ef004076",
          86 => x"13040000",
          87 => x"93040000",
          88 => x"370a00f0",
          89 => x"130b3005",
          90 => x"930ba004",
          91 => x"130c3002",
          92 => x"93092000",
          93 => x"930ca000",
          94 => x"b71a0010",
          95 => x"83274a00",
          96 => x"93c71700",
          97 => x"2322fa00",
          98 => x"ef004053",
          99 => x"1375f50f",
         100 => x"631e6517",
         101 => x"ef008052",
         102 => x"137df50f",
         103 => x"9307fdfc",
         104 => x"93f7f70f",
         105 => x"63e6f910",
         106 => x"93071003",
         107 => x"631afd04",
         108 => x"13052000",
         109 => x"ef004074",
         110 => x"930dd5ff",
         111 => x"13054000",
         112 => x"ef008073",
         113 => x"b70601ff",
         114 => x"b705ffff",
         115 => x"130d0500",
         116 => x"b38dad00",
         117 => x"9386f6ff",
         118 => x"9385f50f",
         119 => x"6398ad05",
         120 => x"130da000",
         121 => x"ef00804d",
         122 => x"1375f50f",
         123 => x"e31ca5ff",
         124 => x"e31604f8",
         125 => x"13850adf",
         126 => x"ef00006c",
         127 => x"6ff01ff8",
         128 => x"93072003",
         129 => x"13052000",
         130 => x"631afd00",
         131 => x"ef00c06e",
         132 => x"930dc5ff",
         133 => x"13056000",
         134 => x"6ff09ffa",
         135 => x"ef00c06d",
         136 => x"930db5ff",
         137 => x"13058000",
         138 => x"6ff09ff9",
         139 => x"1378cdff",
         140 => x"13052000",
         141 => x"2326b100",
         142 => x"2324d100",
         143 => x"23220101",
         144 => x"ef00806b",
         145 => x"03284100",
         146 => x"93070500",
         147 => x"37060001",
         148 => x"13753d00",
         149 => x"03270800",
         150 => x"83268100",
         151 => x"8325c100",
         152 => x"93083000",
         153 => x"1306f6ff",
         154 => x"13031000",
         155 => x"63063503",
         156 => x"630a1503",
         157 => x"630c6500",
         158 => x"137707f0",
         159 => x"b3e7e700",
         160 => x"2320f800",
         161 => x"130d1d00",
         162 => x"6ff05ff5",
         163 => x"3377b700",
         164 => x"93978700",
         165 => x"6ff09ffe",
         166 => x"3377d700",
         167 => x"93970701",
         168 => x"6ff0dffd",
         169 => x"3377c700",
         170 => x"93978701",
         171 => x"6ff01ffd",
         172 => x"93079dfc",
         173 => x"93f7f70f",
         174 => x"63e2f904",
         175 => x"13052000",
         176 => x"ef008063",
         177 => x"93077003",
         178 => x"13058000",
         179 => x"630afd00",
         180 => x"93078003",
         181 => x"13056000",
         182 => x"6304fd00",
         183 => x"13054000",
         184 => x"ef008061",
         185 => x"93040500",
         186 => x"130da000",
         187 => x"ef00003d",
         188 => x"1375f50f",
         189 => x"e31ca5ff",
         190 => x"6ff09fef",
         191 => x"ef00003c",
         192 => x"1375f50f",
         193 => x"e31c95ff",
         194 => x"6ff09fee",
         195 => x"6310750b",
         196 => x"63180400",
         197 => x"37150010",
         198 => x"130505df",
         199 => x"ef00c059",
         200 => x"93050000",
         201 => x"13050000",
         202 => x"ef004054",
         203 => x"b70700f0",
         204 => x"23a20700",
         205 => x"e7800400",
         206 => x"b70700f0",
         207 => x"1307a00a",
         208 => x"23a2e700",
         209 => x"97020000",
         210 => x"93824223",
         211 => x"73905230",
         212 => x"b7190010",
         213 => x"130589dd",
         214 => x"ef000056",
         215 => x"13040000",
         216 => x"371b0010",
         217 => x"b71b0010",
         218 => x"938959c9",
         219 => x"b7170010",
         220 => x"138547df",
         221 => x"ef004054",
         222 => x"93059002",
         223 => x"13054101",
         224 => x"ef00c035",
         225 => x"b7170010",
         226 => x"130a0500",
         227 => x"938587df",
         228 => x"13054101",
         229 => x"ef00802f",
         230 => x"631e0500",
         231 => x"37150010",
         232 => x"1305c5df",
         233 => x"ef004051",
         234 => x"6f00c003",
         235 => x"e31285e5",
         236 => x"6ff09ff8",
         237 => x"b7170010",
         238 => x"938587ee",
         239 => x"13054101",
         240 => x"ef00c02c",
         241 => x"63140502",
         242 => x"93050000",
         243 => x"ef00004a",
         244 => x"b70700f0",
         245 => x"23a20700",
         246 => x"93020000",
         247 => x"73905230",
         248 => x"e7800400",
         249 => x"e3040af8",
         250 => x"6f004018",
         251 => x"b7170010",
         252 => x"13063000",
         253 => x"9385c7ee",
         254 => x"13054101",
         255 => x"ef001001",
         256 => x"63100504",
         257 => x"93050000",
         258 => x"13057101",
         259 => x"ef00005b",
         260 => x"93773500",
         261 => x"13040500",
         262 => x"63940706",
         263 => x"93058000",
         264 => x"ef00406e",
         265 => x"37150010",
         266 => x"130505ef",
         267 => x"ef00c048",
         268 => x"03250400",
         269 => x"93058000",
         270 => x"ef00c06c",
         271 => x"6ff09ffa",
         272 => x"13063000",
         273 => x"9305cbf0",
         274 => x"13054101",
         275 => x"ef00007c",
         276 => x"631e0502",
         277 => x"93050101",
         278 => x"13057101",
         279 => x"ef000056",
         280 => x"93773500",
         281 => x"13040500",
         282 => x"639c0700",
         283 => x"03250101",
         284 => x"93050000",
         285 => x"ef008054",
         286 => x"2320a400",
         287 => x"6ff09ff6",
         288 => x"37150010",
         289 => x"130545ef",
         290 => x"6ff0dff1",
         291 => x"13063000",
         292 => x"93850bf1",
         293 => x"13054101",
         294 => x"ef004077",
         295 => x"83474101",
         296 => x"1307e006",
         297 => x"630c0508",
         298 => x"639ae70a",
         299 => x"93773400",
         300 => x"e39807fc",
         301 => x"130c0404",
         302 => x"b71c0010",
         303 => x"371d0010",
         304 => x"930d80ff",
         305 => x"93058000",
         306 => x"13050400",
         307 => x"ef008063",
         308 => x"13850cef",
         309 => x"ef00403e",
         310 => x"83270400",
         311 => x"93058000",
         312 => x"130a8001",
         313 => x"13850700",
         314 => x"2322f100",
         315 => x"ef008061",
         316 => x"13054df1",
         317 => x"ef00403c",
         318 => x"b70a00ff",
         319 => x"83274100",
         320 => x"33f55701",
         321 => x"33554501",
         322 => x"b3063501",
         323 => x"83c60600",
         324 => x"93f67609",
         325 => x"63800604",
         326 => x"130a8aff",
         327 => x"ef00c037",
         328 => x"93da8a00",
         329 => x"e31cbafd",
         330 => x"13044400",
         331 => x"130589dd",
         332 => x"ef008038",
         333 => x"e3188cf8",
         334 => x"6ff05fe3",
         335 => x"e388e7f6",
         336 => x"93050000",
         337 => x"13057101",
         338 => x"ef004047",
         339 => x"13040500",
         340 => x"6ff0dff5",
         341 => x"1305e002",
         342 => x"6ff01ffc",
         343 => x"e3080ae0",
         344 => x"37150010",
         345 => x"130585f1",
         346 => x"ef000035",
         347 => x"130589dd",
         348 => x"ef008034",
         349 => x"6ff09fdf",
         350 => x"130101fb",
         351 => x"23261104",
         352 => x"23245104",
         353 => x"23226104",
         354 => x"23207104",
         355 => x"232e8102",
         356 => x"232c9102",
         357 => x"232aa102",
         358 => x"2328b102",
         359 => x"2326c102",
         360 => x"2324d102",
         361 => x"2322e102",
         362 => x"2320f102",
         363 => x"232e0101",
         364 => x"232c1101",
         365 => x"232ac101",
         366 => x"2328d101",
         367 => x"2326e101",
         368 => x"2324f101",
         369 => x"73241034",
         370 => x"f3242034",
         371 => x"37150010",
         372 => x"130545da",
         373 => x"ef00402e",
         374 => x"93058000",
         375 => x"13850400",
         376 => x"ef004052",
         377 => x"37150010",
         378 => x"130585dd",
         379 => x"ef00c02c",
         380 => x"13044400",
         381 => x"73101434",
         382 => x"0324c103",
         383 => x"8320c104",
         384 => x"83228104",
         385 => x"03234104",
         386 => x"83230104",
         387 => x"83248103",
         388 => x"03254103",
         389 => x"83250103",
         390 => x"0326c102",
         391 => x"83268102",
         392 => x"03274102",
         393 => x"83270102",
         394 => x"0328c101",
         395 => x"83288101",
         396 => x"032e4101",
         397 => x"832e0101",
         398 => x"032fc100",
         399 => x"832f8100",
         400 => x"13010105",
         401 => x"73002030",
         402 => x"6f000000",
         403 => x"13030500",
         404 => x"630a0600",
         405 => x"2300b300",
         406 => x"1306f6ff",
         407 => x"13031300",
         408 => x"e31a06fe",
         409 => x"67800000",
         410 => x"13030500",
         411 => x"630e0600",
         412 => x"83830500",
         413 => x"23007300",
         414 => x"1306f6ff",
         415 => x"13031300",
         416 => x"93851500",
         417 => x"e31606fe",
         418 => x"67800000",
         419 => x"03460500",
         420 => x"83c60500",
         421 => x"13051500",
         422 => x"93851500",
         423 => x"6314d600",
         424 => x"e31606fe",
         425 => x"3305d640",
         426 => x"67800000",
         427 => x"b70700f0",
         428 => x"03a54702",
         429 => x"13758500",
         430 => x"67800000",
         431 => x"370700f0",
         432 => x"13070702",
         433 => x"83274700",
         434 => x"93f78700",
         435 => x"e38c07fe",
         436 => x"03258700",
         437 => x"1375f50f",
         438 => x"67800000",
         439 => x"130101fd",
         440 => x"232e3101",
         441 => x"b7190010",
         442 => x"23248102",
         443 => x"23229102",
         444 => x"23202103",
         445 => x"232c4101",
         446 => x"232a5101",
         447 => x"23286101",
         448 => x"23267101",
         449 => x"23261102",
         450 => x"93040500",
         451 => x"13040000",
         452 => x"938989c4",
         453 => x"13095001",
         454 => x"138bf5ff",
         455 => x"130a2000",
         456 => x"930a2001",
         457 => x"b71b0010",
         458 => x"eff05ff9",
         459 => x"1377f50f",
         460 => x"6340e902",
         461 => x"6352ea02",
         462 => x"9307d7ff",
         463 => x"63eefa00",
         464 => x"93972700",
         465 => x"b387f900",
         466 => x"83a70700",
         467 => x"67800700",
         468 => x"9307f007",
         469 => x"630cf706",
         470 => x"6352640f",
         471 => x"9377f50f",
         472 => x"938607fe",
         473 => x"93f6f60f",
         474 => x"1306e005",
         475 => x"e36ed6fa",
         476 => x"b3868400",
         477 => x"2380f600",
         478 => x"13050700",
         479 => x"13041400",
         480 => x"ef008011",
         481 => x"6ff05ffa",
         482 => x"b3848400",
         483 => x"37150010",
         484 => x"23800400",
         485 => x"130585dd",
         486 => x"ef000012",
         487 => x"8320c102",
         488 => x"13050400",
         489 => x"03248102",
         490 => x"83244102",
         491 => x"03290102",
         492 => x"8329c101",
         493 => x"032a8101",
         494 => x"832a4101",
         495 => x"032b0101",
         496 => x"832bc100",
         497 => x"13010103",
         498 => x"67800000",
         499 => x"635a8002",
         500 => x"1305f007",
         501 => x"ef00400c",
         502 => x"1304f4ff",
         503 => x"6ff0dff4",
         504 => x"13858bd9",
         505 => x"ef00400d",
         506 => x"eff05fed",
         507 => x"1377f50f",
         508 => x"13040000",
         509 => x"e350e9f4",
         510 => x"9307f007",
         511 => x"e31ef7f4",
         512 => x"23248101",
         513 => x"130c5001",
         514 => x"13057000",
         515 => x"ef00c008",
         516 => x"eff0dfea",
         517 => x"1377f50f",
         518 => x"6348ec02",
         519 => x"032c8100",
         520 => x"6ff05ff1",
         521 => x"635a8002",
         522 => x"1305f007",
         523 => x"1304f4ff",
         524 => x"ef008006",
         525 => x"e31a04fe",
         526 => x"6ff01fef",
         527 => x"13057000",
         528 => x"ef008005",
         529 => x"6ff05fee",
         530 => x"9307f007",
         531 => x"e30ef7fa",
         532 => x"032c8100",
         533 => x"6ff05ff0",
         534 => x"eff05fe6",
         535 => x"1377f50f",
         536 => x"93075001",
         537 => x"e3d8e7ec",
         538 => x"6ff01ff9",
         539 => x"f32710fc",
         540 => x"63960700",
         541 => x"b7f7fa02",
         542 => x"93870708",
         543 => x"63060500",
         544 => x"33d5a702",
         545 => x"1305f5ff",
         546 => x"b70700f0",
         547 => x"23a6a702",
         548 => x"23a0b702",
         549 => x"67800000",
         550 => x"370700f0",
         551 => x"1375f50f",
         552 => x"13070702",
         553 => x"2324a700",
         554 => x"83274700",
         555 => x"93f70701",
         556 => x"e38c07fe",
         557 => x"67800000",
         558 => x"630e0502",
         559 => x"130101ff",
         560 => x"23248100",
         561 => x"23261100",
         562 => x"13040500",
         563 => x"03450500",
         564 => x"630a0500",
         565 => x"13041400",
         566 => x"eff01ffc",
         567 => x"03450400",
         568 => x"e31a05fe",
         569 => x"8320c100",
         570 => x"03248100",
         571 => x"13010101",
         572 => x"67800000",
         573 => x"67800000",
         574 => x"130101fe",
         575 => x"232e1100",
         576 => x"232c8100",
         577 => x"6350a00a",
         578 => x"23263101",
         579 => x"b7190010",
         580 => x"232a9100",
         581 => x"23282101",
         582 => x"23244101",
         583 => x"13090500",
         584 => x"93040000",
         585 => x"13040000",
         586 => x"938959c9",
         587 => x"130a1000",
         588 => x"6f000001",
         589 => x"3364c400",
         590 => x"93841400",
         591 => x"63029904",
         592 => x"eff0dfd7",
         593 => x"b387a900",
         594 => x"83c70700",
         595 => x"130605fd",
         596 => x"13144400",
         597 => x"13f74700",
         598 => x"93f64704",
         599 => x"e31c07fc",
         600 => x"93f73700",
         601 => x"e38a06fc",
         602 => x"63944701",
         603 => x"13050502",
         604 => x"130595fa",
         605 => x"93841400",
         606 => x"3364a400",
         607 => x"e31299fc",
         608 => x"8320c101",
         609 => x"13050400",
         610 => x"03248101",
         611 => x"83244101",
         612 => x"03290101",
         613 => x"8329c100",
         614 => x"032a8100",
         615 => x"13010102",
         616 => x"67800000",
         617 => x"13040000",
         618 => x"8320c101",
         619 => x"13050400",
         620 => x"03248101",
         621 => x"13010102",
         622 => x"67800000",
         623 => x"83470500",
         624 => x"37160010",
         625 => x"130656c9",
         626 => x"3307f600",
         627 => x"03470700",
         628 => x"93060500",
         629 => x"13758700",
         630 => x"630e0500",
         631 => x"83c71600",
         632 => x"93861600",
         633 => x"3307f600",
         634 => x"03470700",
         635 => x"13758700",
         636 => x"e31605fe",
         637 => x"13754704",
         638 => x"630a0506",
         639 => x"13050000",
         640 => x"13031000",
         641 => x"6f000002",
         642 => x"83c71600",
         643 => x"33e5a800",
         644 => x"93861600",
         645 => x"3307f600",
         646 => x"03470700",
         647 => x"13784704",
         648 => x"63000804",
         649 => x"13784700",
         650 => x"938807fd",
         651 => x"13773700",
         652 => x"13154500",
         653 => x"e31a08fc",
         654 => x"63146700",
         655 => x"93870702",
         656 => x"938797fa",
         657 => x"33e5a700",
         658 => x"83c71600",
         659 => x"93861600",
         660 => x"3307f600",
         661 => x"03470700",
         662 => x"13784704",
         663 => x"e31408fc",
         664 => x"63840500",
         665 => x"23a0d500",
         666 => x"67800000",
         667 => x"13050000",
         668 => x"6ff01fff",
         669 => x"130101fe",
         670 => x"232e1100",
         671 => x"23220100",
         672 => x"23240100",
         673 => x"23260100",
         674 => x"63040506",
         675 => x"232c8100",
         676 => x"93070500",
         677 => x"13040500",
         678 => x"63440504",
         679 => x"13074100",
         680 => x"1306a000",
         681 => x"13089000",
         682 => x"b3f6c702",
         683 => x"13050700",
         684 => x"1307f7ff",
         685 => x"93850700",
         686 => x"93860603",
         687 => x"a305d700",
         688 => x"b3d7c702",
         689 => x"e362b8fe",
         690 => x"3305c500",
         691 => x"eff0dfde",
         692 => x"8320c101",
         693 => x"03248101",
         694 => x"13010102",
         695 => x"67800000",
         696 => x"1305d002",
         697 => x"eff05fdb",
         698 => x"b3078040",
         699 => x"6ff01ffb",
         700 => x"13050003",
         701 => x"eff05fda",
         702 => x"8320c101",
         703 => x"13010102",
         704 => x"67800000",
         705 => x"130101fe",
         706 => x"232e1100",
         707 => x"23220100",
         708 => x"23240100",
         709 => x"23060100",
         710 => x"9387f5ff",
         711 => x"13077000",
         712 => x"6376f700",
         713 => x"93077000",
         714 => x"93058000",
         715 => x"13074100",
         716 => x"b307f700",
         717 => x"b385b740",
         718 => x"13069003",
         719 => x"9376f500",
         720 => x"13870603",
         721 => x"6374e600",
         722 => x"13877605",
         723 => x"2380e700",
         724 => x"9387f7ff",
         725 => x"13554500",
         726 => x"e392f5fe",
         727 => x"13054100",
         728 => x"eff09fd5",
         729 => x"8320c101",
         730 => x"13010102",
         731 => x"67800000",
         732 => x"130101ff",
         733 => x"23248100",
         734 => x"23229100",
         735 => x"37140010",
         736 => x"b7140010",
         737 => x"9387c4f1",
         738 => x"1304c4f1",
         739 => x"3304f440",
         740 => x"23202101",
         741 => x"23261100",
         742 => x"13542440",
         743 => x"9384c4f1",
         744 => x"13090000",
         745 => x"63108904",
         746 => x"b7140010",
         747 => x"37140010",
         748 => x"9387c4f1",
         749 => x"1304c4f1",
         750 => x"3304f440",
         751 => x"13542440",
         752 => x"9384c4f1",
         753 => x"13090000",
         754 => x"63188902",
         755 => x"8320c100",
         756 => x"03248100",
         757 => x"83244100",
         758 => x"03290100",
         759 => x"13010101",
         760 => x"67800000",
         761 => x"83a70400",
         762 => x"13091900",
         763 => x"93844400",
         764 => x"e7800700",
         765 => x"6ff01ffb",
         766 => x"83a70400",
         767 => x"13091900",
         768 => x"93844400",
         769 => x"e7800700",
         770 => x"6ff01ffc",
         771 => x"630a0602",
         772 => x"1306f6ff",
         773 => x"13070000",
         774 => x"b307e500",
         775 => x"b386e500",
         776 => x"83c70700",
         777 => x"83c60600",
         778 => x"6398d700",
         779 => x"6306c700",
         780 => x"13071700",
         781 => x"e39207fe",
         782 => x"3385d740",
         783 => x"67800000",
         784 => x"13050000",
         785 => x"67800000",
         786 => x"e0070010",
         787 => x"58070010",
         788 => x"58070010",
         789 => x"58070010",
         790 => x"58070010",
         791 => x"cc070010",
         792 => x"58070010",
         793 => x"88070010",
         794 => x"58070010",
         795 => x"58070010",
         796 => x"88070010",
         797 => x"58070010",
         798 => x"58070010",
         799 => x"58070010",
         800 => x"58070010",
         801 => x"58070010",
         802 => x"58070010",
         803 => x"58070010",
         804 => x"24080010",
         805 => x"00202020",
         806 => x"20202020",
         807 => x"20202828",
         808 => x"28282820",
         809 => x"20202020",
         810 => x"20202020",
         811 => x"20202020",
         812 => x"20202020",
         813 => x"20881010",
         814 => x"10101010",
         815 => x"10101010",
         816 => x"10101010",
         817 => x"10040404",
         818 => x"04040404",
         819 => x"04040410",
         820 => x"10101010",
         821 => x"10104141",
         822 => x"41414141",
         823 => x"01010101",
         824 => x"01010101",
         825 => x"01010101",
         826 => x"01010101",
         827 => x"01010101",
         828 => x"10101010",
         829 => x"10104242",
         830 => x"42424242",
         831 => x"02020202",
         832 => x"02020202",
         833 => x"02020202",
         834 => x"02020202",
         835 => x"02020202",
         836 => x"10101010",
         837 => x"20000000",
         838 => x"00000000",
         839 => x"00000000",
         840 => x"00000000",
         841 => x"00000000",
         842 => x"00000000",
         843 => x"00000000",
         844 => x"00000000",
         845 => x"00000000",
         846 => x"00000000",
         847 => x"00000000",
         848 => x"00000000",
         849 => x"00000000",
         850 => x"00000000",
         851 => x"00000000",
         852 => x"00000000",
         853 => x"00000000",
         854 => x"00000000",
         855 => x"00000000",
         856 => x"00000000",
         857 => x"00000000",
         858 => x"00000000",
         859 => x"00000000",
         860 => x"00000000",
         861 => x"00000000",
         862 => x"00000000",
         863 => x"00000000",
         864 => x"00000000",
         865 => x"00000000",
         866 => x"00000000",
         867 => x"00000000",
         868 => x"00000000",
         869 => x"00000000",
         870 => x"3c627265",
         871 => x"616b3e0d",
         872 => x"0a000000",
         873 => x"54726170",
         874 => x"3a206d63",
         875 => x"61757365",
         876 => x"203d2030",
         877 => x"78000000",
         878 => x"0d0a5448",
         879 => x"55415320",
         880 => x"52495343",
         881 => x"2d562042",
         882 => x"6f6f746c",
         883 => x"6f616465",
         884 => x"72207630",
         885 => x"2e362e31",
         886 => x"0d0a0000",
         887 => x"436c6f63",
         888 => x"6b206672",
         889 => x"65717565",
         890 => x"6e63793a",
         891 => x"20000000",
         892 => x"3f0a0000",
         893 => x"3e200000",
         894 => x"68000000",
         895 => x"48656c70",
         896 => x"3a0d0a20",
         897 => x"68202020",
         898 => x"20202020",
         899 => x"20202020",
         900 => x"20202020",
         901 => x"202d2074",
         902 => x"68697320",
         903 => x"68656c70",
         904 => x"0d0a2072",
         905 => x"20202020",
         906 => x"20202020",
         907 => x"20202020",
         908 => x"20202020",
         909 => x"2d207275",
         910 => x"6e206170",
         911 => x"706c6963",
         912 => x"6174696f",
         913 => x"6e0d0a20",
         914 => x"7277203c",
         915 => x"61646472",
         916 => x"3e202020",
         917 => x"20202020",
         918 => x"202d2072",
         919 => x"65616420",
         920 => x"776f7264",
         921 => x"2066726f",
         922 => x"6d206164",
         923 => x"64720d0a",
         924 => x"20777720",
         925 => x"3c616464",
         926 => x"723e203c",
         927 => x"64617461",
         928 => x"3e202d20",
         929 => x"77726974",
         930 => x"6520776f",
         931 => x"72642064",
         932 => x"61746120",
         933 => x"61742061",
         934 => x"6464720d",
         935 => x"0a206477",
         936 => x"203c6164",
         937 => x"64723e20",
         938 => x"20202020",
         939 => x"2020202d",
         940 => x"2064756d",
         941 => x"70203136",
         942 => x"20776f72",
         943 => x"64730d0a",
         944 => x"206e2020",
         945 => x"20202020",
         946 => x"20202020",
         947 => x"20202020",
         948 => x"20202d20",
         949 => x"64756d70",
         950 => x"206e6578",
         951 => x"74203136",
         952 => x"20776f72",
         953 => x"64730000",
         954 => x"72000000",
         955 => x"72772000",
         956 => x"3a200000",
         957 => x"4e6f7420",
         958 => x"6f6e2034",
         959 => x"2d627974",
         960 => x"6520626f",
         961 => x"756e6461",
         962 => x"72792100",
         963 => x"77772000",
         964 => x"64772000",
         965 => x"20200000",
         966 => x"3f3f0000",
         967 => x"00000000"
            );
end package bootrom_image;
