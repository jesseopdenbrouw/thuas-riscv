-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Tue Nov  7 10:56:02 2023


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382422d",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"13868187",
           8 => x"9387819c",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13858187",
          13 => x"ef10c032",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93878187",
          17 => x"637cf600",
          18 => x"b7450000",
          19 => x"3386c740",
          20 => x"9385c5be",
          21 => x"13050500",
          22 => x"ef104032",
          23 => x"ef20402e",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef100070",
          29 => x"ef10d027",
          30 => x"6f10c064",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef10c068",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"232c4101",
          40 => x"130a0500",
          41 => x"37450000",
          42 => x"130585a3",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"13044100",
          50 => x"ef108066",
          51 => x"37390000",
          52 => x"9309c1ff",
          53 => x"93070400",
          54 => x"1309c97c",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef100063",
          65 => x"37450000",
          66 => x"1305c5a4",
          67 => x"ef104062",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef10c05f",
          78 => x"37450000",
          79 => x"130585a5",
          80 => x"ef10005f",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74708",
          91 => x"b70600f0",
          92 => x"1377f7fe",
          93 => x"23a2e708",
          94 => x"83a74600",
          95 => x"93c71700",
          96 => x"23a2f600",
          97 => x"67800000",
          98 => x"370700f0",
          99 => x"83274700",
         100 => x"93e70720",
         101 => x"2322f700",
         102 => x"6f000000",
         103 => x"b70700f0",
         104 => x"b70500f0",
         105 => x"370500f0",
         106 => x"9387470f",
         107 => x"9385050f",
         108 => x"83a60700",
         109 => x"03a60500",
         110 => x"03a70700",
         111 => x"e31ad7fe",
         112 => x"b7870100",
         113 => x"b70500f0",
         114 => x"1308f0ff",
         115 => x"9387076a",
         116 => x"23ae050f",
         117 => x"b307f600",
         118 => x"b70600f0",
         119 => x"23ac060f",
         120 => x"33b6c700",
         121 => x"23acf60e",
         122 => x"3306e600",
         123 => x"23aec50e",
         124 => x"83274500",
         125 => x"93c72700",
         126 => x"2322f500",
         127 => x"67800000",
         128 => x"b70700f0",
         129 => x"03a74702",
         130 => x"b70600f0",
         131 => x"93870702",
         132 => x"13770701",
         133 => x"630a0700",
         134 => x"03a74600",
         135 => x"13478700",
         136 => x"23a2e600",
         137 => x"83a78700",
         138 => x"67800000",
         139 => x"b70700f0",
         140 => x"03a7470a",
         141 => x"b70600f0",
         142 => x"1377f7f0",
         143 => x"23a2e70a",
         144 => x"83a74600",
         145 => x"93c74700",
         146 => x"23a2f600",
         147 => x"67800000",
         148 => x"b70700f0",
         149 => x"03a74706",
         150 => x"b70600f0",
         151 => x"137777ff",
         152 => x"23a2e706",
         153 => x"83a74600",
         154 => x"93c70701",
         155 => x"23a2f600",
         156 => x"67800000",
         157 => x"b70700f0",
         158 => x"03a74704",
         159 => x"b70600f0",
         160 => x"137777ff",
         161 => x"23a2e704",
         162 => x"83a74600",
         163 => x"93c70702",
         164 => x"23a2f600",
         165 => x"67800000",
         166 => x"b70700f0",
         167 => x"03a74705",
         168 => x"b70600f0",
         169 => x"137777ff",
         170 => x"23aae704",
         171 => x"83a74600",
         172 => x"93c70708",
         173 => x"23a2f600",
         174 => x"67800000",
         175 => x"b70700f0",
         176 => x"23ae0700",
         177 => x"03a74700",
         178 => x"13470704",
         179 => x"23a2e700",
         180 => x"67800000",
         181 => x"6f000000",
         182 => x"13050000",
         183 => x"67800000",
         184 => x"13050000",
         185 => x"67800000",
         186 => x"130101f7",
         187 => x"23221100",
         188 => x"23242100",
         189 => x"23263100",
         190 => x"23284100",
         191 => x"232a5100",
         192 => x"232c6100",
         193 => x"232e7100",
         194 => x"23208102",
         195 => x"23229102",
         196 => x"2324a102",
         197 => x"2326b102",
         198 => x"2328c102",
         199 => x"232ad102",
         200 => x"232ce102",
         201 => x"232ef102",
         202 => x"23200105",
         203 => x"23221105",
         204 => x"23242105",
         205 => x"23263105",
         206 => x"23284105",
         207 => x"232a5105",
         208 => x"232c6105",
         209 => x"232e7105",
         210 => x"23208107",
         211 => x"23229107",
         212 => x"2324a107",
         213 => x"2326b107",
         214 => x"2328c107",
         215 => x"232ad107",
         216 => x"232ce107",
         217 => x"232ef107",
         218 => x"f3222034",
         219 => x"23205108",
         220 => x"f3221034",
         221 => x"23225108",
         222 => x"83a20200",
         223 => x"23245108",
         224 => x"f3223034",
         225 => x"23265108",
         226 => x"f3272034",
         227 => x"1307b000",
         228 => x"6374f70c",
         229 => x"37070080",
         230 => x"130797ff",
         231 => x"b387e700",
         232 => x"13074001",
         233 => x"636ef700",
         234 => x"37370000",
         235 => x"93972700",
         236 => x"1307077e",
         237 => x"b387e700",
         238 => x"83a70700",
         239 => x"67800700",
         240 => x"03258102",
         241 => x"83220108",
         242 => x"63c80200",
         243 => x"f3221034",
         244 => x"93824200",
         245 => x"73901234",
         246 => x"832fc107",
         247 => x"032f8107",
         248 => x"832e4107",
         249 => x"032e0107",
         250 => x"832dc106",
         251 => x"032d8106",
         252 => x"832c4106",
         253 => x"032c0106",
         254 => x"832bc105",
         255 => x"032b8105",
         256 => x"832a4105",
         257 => x"032a0105",
         258 => x"8329c104",
         259 => x"03298104",
         260 => x"83284104",
         261 => x"03280104",
         262 => x"8327c103",
         263 => x"03278103",
         264 => x"83264103",
         265 => x"03260103",
         266 => x"8325c102",
         267 => x"83244102",
         268 => x"03240102",
         269 => x"8323c101",
         270 => x"03238101",
         271 => x"83224101",
         272 => x"03220101",
         273 => x"8321c100",
         274 => x"03218100",
         275 => x"83204100",
         276 => x"13010109",
         277 => x"73002030",
         278 => x"93061000",
         279 => x"e3f2f6f6",
         280 => x"e360f7f6",
         281 => x"37470000",
         282 => x"93972700",
         283 => x"13074783",
         284 => x"b387e700",
         285 => x"83a70700",
         286 => x"67800700",
         287 => x"eff05fdd",
         288 => x"03258102",
         289 => x"6ff01ff4",
         290 => x"eff05fd1",
         291 => x"03258102",
         292 => x"6ff05ff3",
         293 => x"eff09fe2",
         294 => x"03258102",
         295 => x"6ff09ff2",
         296 => x"eff05fcc",
         297 => x"03258102",
         298 => x"6ff0dff1",
         299 => x"eff01fd8",
         300 => x"03258102",
         301 => x"6ff01ff1",
         302 => x"eff09fd4",
         303 => x"03258102",
         304 => x"6ff05ff0",
         305 => x"eff05fdd",
         306 => x"03258102",
         307 => x"6ff09fef",
         308 => x"eff05fda",
         309 => x"03258102",
         310 => x"6ff0dfee",
         311 => x"13050100",
         312 => x"eff09fbb",
         313 => x"03258102",
         314 => x"6ff0dfed",
         315 => x"9307900a",
         316 => x"6380f814",
         317 => x"63d81703",
         318 => x"9307600d",
         319 => x"638ef818",
         320 => x"938808c0",
         321 => x"9307f000",
         322 => x"63e01705",
         323 => x"b7470000",
         324 => x"93874786",
         325 => x"93982800",
         326 => x"b388f800",
         327 => x"83a70800",
         328 => x"67800700",
         329 => x"938878fc",
         330 => x"93074002",
         331 => x"63ee1701",
         332 => x"b7470000",
         333 => x"9387478a",
         334 => x"93982800",
         335 => x"b388f800",
         336 => x"83a70800",
         337 => x"67800700",
         338 => x"ef10105f",
         339 => x"93078005",
         340 => x"2320f500",
         341 => x"9307f0ff",
         342 => x"13850700",
         343 => x"6ff09fe6",
         344 => x"b7270000",
         345 => x"23a2f500",
         346 => x"93070000",
         347 => x"13850700",
         348 => x"6ff05fe5",
         349 => x"93070000",
         350 => x"13850700",
         351 => x"6ff09fe4",
         352 => x"ef10905b",
         353 => x"93079000",
         354 => x"2320f500",
         355 => x"9307f0ff",
         356 => x"13850700",
         357 => x"6ff01fe3",
         358 => x"ef10105a",
         359 => x"9307f001",
         360 => x"2320f500",
         361 => x"9307f0ff",
         362 => x"13850700",
         363 => x"6ff09fe1",
         364 => x"ef109058",
         365 => x"9307d000",
         366 => x"2320f500",
         367 => x"9307f0ff",
         368 => x"13850700",
         369 => x"6ff01fe0",
         370 => x"ef101057",
         371 => x"93072000",
         372 => x"2320f500",
         373 => x"9307f0ff",
         374 => x"13850700",
         375 => x"6ff09fde",
         376 => x"13090600",
         377 => x"13840500",
         378 => x"635cc000",
         379 => x"b384c500",
         380 => x"eff09fa8",
         381 => x"2300a400",
         382 => x"13041400",
         383 => x"e39a84fe",
         384 => x"13050900",
         385 => x"6ff01fdc",
         386 => x"13090600",
         387 => x"13840500",
         388 => x"e358c0fe",
         389 => x"b384c500",
         390 => x"03450400",
         391 => x"13041400",
         392 => x"eff0dfa5",
         393 => x"e39a84fe",
         394 => x"13050900",
         395 => x"6ff09fd9",
         396 => x"13090000",
         397 => x"93040500",
         398 => x"13040900",
         399 => x"93090900",
         400 => x"93070900",
         401 => x"732410c8",
         402 => x"f32910c0",
         403 => x"f32710c8",
         404 => x"e31af4fe",
         405 => x"37460f00",
         406 => x"13060624",
         407 => x"93060000",
         408 => x"13850900",
         409 => x"93050400",
         410 => x"ef005011",
         411 => x"37460f00",
         412 => x"23a4a400",
         413 => x"13060624",
         414 => x"93060000",
         415 => x"13850900",
         416 => x"93050400",
         417 => x"ef00804c",
         418 => x"23a0a400",
         419 => x"23a2b400",
         420 => x"13050900",
         421 => x"6ff01fd3",
         422 => x"63180500",
         423 => x"1385819c",
         424 => x"13050500",
         425 => x"6ff01fd2",
         426 => x"b7870020",
         427 => x"93870700",
         428 => x"13070040",
         429 => x"b387e740",
         430 => x"e364f5fe",
         431 => x"ef10d047",
         432 => x"9307c000",
         433 => x"2320f500",
         434 => x"1305f0ff",
         435 => x"13050500",
         436 => x"6ff05fcf",
         437 => x"13030500",
         438 => x"138e0500",
         439 => x"93080000",
         440 => x"63dc0500",
         441 => x"b337a000",
         442 => x"330eb040",
         443 => x"330efe40",
         444 => x"3303a040",
         445 => x"9308f0ff",
         446 => x"63dc0600",
         447 => x"b337c000",
         448 => x"b306d040",
         449 => x"93c8f8ff",
         450 => x"b386f640",
         451 => x"3306c040",
         452 => x"13070600",
         453 => x"13080300",
         454 => x"93070e00",
         455 => x"639c0628",
         456 => x"b7450000",
         457 => x"93858593",
         458 => x"6376ce0e",
         459 => x"b7060100",
         460 => x"6378d60c",
         461 => x"93360610",
         462 => x"93b61600",
         463 => x"93963600",
         464 => x"3355d600",
         465 => x"b385a500",
         466 => x"83c50500",
         467 => x"13050002",
         468 => x"b386d500",
         469 => x"b305d540",
         470 => x"630cd500",
         471 => x"b317be00",
         472 => x"b356d300",
         473 => x"3317b600",
         474 => x"b3e7f600",
         475 => x"3318b300",
         476 => x"93550701",
         477 => x"33deb702",
         478 => x"13160701",
         479 => x"13560601",
         480 => x"b3f7b702",
         481 => x"13050e00",
         482 => x"3303c603",
         483 => x"93960701",
         484 => x"93570801",
         485 => x"b3e7d700",
         486 => x"63fe6700",
         487 => x"b307f700",
         488 => x"1305feff",
         489 => x"63e8e700",
         490 => x"63f66700",
         491 => x"1305eeff",
         492 => x"b387e700",
         493 => x"b3876740",
         494 => x"33d3b702",
         495 => x"13180801",
         496 => x"13580801",
         497 => x"b3f7b702",
         498 => x"b3066602",
         499 => x"93970701",
         500 => x"3368f800",
         501 => x"93070300",
         502 => x"637cd800",
         503 => x"33080701",
         504 => x"9307f3ff",
         505 => x"6366e800",
         506 => x"6374d800",
         507 => x"9307e3ff",
         508 => x"13150501",
         509 => x"3365f500",
         510 => x"93050000",
         511 => x"6f00000e",
         512 => x"37050001",
         513 => x"93068001",
         514 => x"e37ca6f2",
         515 => x"93060001",
         516 => x"6ff01ff3",
         517 => x"93060000",
         518 => x"630c0600",
         519 => x"b7070100",
         520 => x"637af60c",
         521 => x"93360610",
         522 => x"93b61600",
         523 => x"93963600",
         524 => x"b357d600",
         525 => x"b385f500",
         526 => x"83c70500",
         527 => x"b387d700",
         528 => x"93060002",
         529 => x"b385f640",
         530 => x"6390f60c",
         531 => x"b307ce40",
         532 => x"93051000",
         533 => x"13530701",
         534 => x"b3de6702",
         535 => x"13160701",
         536 => x"13560601",
         537 => x"93560801",
         538 => x"b3f76702",
         539 => x"13850e00",
         540 => x"330ed603",
         541 => x"93970701",
         542 => x"b3e7f600",
         543 => x"63fec701",
         544 => x"b307f700",
         545 => x"1385feff",
         546 => x"63e8e700",
         547 => x"63f6c701",
         548 => x"1385eeff",
         549 => x"b387e700",
         550 => x"b387c741",
         551 => x"33de6702",
         552 => x"13180801",
         553 => x"13580801",
         554 => x"b3f76702",
         555 => x"b306c603",
         556 => x"93970701",
         557 => x"3368f800",
         558 => x"93070e00",
         559 => x"637cd800",
         560 => x"33080701",
         561 => x"9307feff",
         562 => x"6366e800",
         563 => x"6374d800",
         564 => x"9307eeff",
         565 => x"13150501",
         566 => x"3365f500",
         567 => x"638a0800",
         568 => x"b337a000",
         569 => x"b305b040",
         570 => x"b385f540",
         571 => x"3305a040",
         572 => x"67800000",
         573 => x"b7070001",
         574 => x"93068001",
         575 => x"e37af6f2",
         576 => x"93060001",
         577 => x"6ff0dff2",
         578 => x"3317b600",
         579 => x"b356fe00",
         580 => x"13550701",
         581 => x"331ebe00",
         582 => x"b357f300",
         583 => x"b3e7c701",
         584 => x"33dea602",
         585 => x"13160701",
         586 => x"13560601",
         587 => x"3318b300",
         588 => x"b3f6a602",
         589 => x"3303c603",
         590 => x"93950601",
         591 => x"93d60701",
         592 => x"b3e6b600",
         593 => x"93050e00",
         594 => x"63fe6600",
         595 => x"b306d700",
         596 => x"9305feff",
         597 => x"63e8e600",
         598 => x"63f66600",
         599 => x"9305eeff",
         600 => x"b386e600",
         601 => x"b3866640",
         602 => x"33d3a602",
         603 => x"93970701",
         604 => x"93d70701",
         605 => x"b3f6a602",
         606 => x"33066602",
         607 => x"93960601",
         608 => x"b3e7d700",
         609 => x"93060300",
         610 => x"63fec700",
         611 => x"b307f700",
         612 => x"9306f3ff",
         613 => x"63e8e700",
         614 => x"63f6c700",
         615 => x"9306e3ff",
         616 => x"b387e700",
         617 => x"93950501",
         618 => x"b387c740",
         619 => x"b3e5d500",
         620 => x"6ff05fea",
         621 => x"6366de18",
         622 => x"b7070100",
         623 => x"63f4f604",
         624 => x"13b70610",
         625 => x"13371700",
         626 => x"13173700",
         627 => x"b7470000",
         628 => x"b3d5e600",
         629 => x"93878793",
         630 => x"b387b700",
         631 => x"83c70700",
         632 => x"b387e700",
         633 => x"13070002",
         634 => x"b305f740",
         635 => x"6316f702",
         636 => x"13051000",
         637 => x"e3e4c6ef",
         638 => x"3335c300",
         639 => x"13351500",
         640 => x"6ff0dfed",
         641 => x"b7070001",
         642 => x"13078001",
         643 => x"e3f0f6fc",
         644 => x"13070001",
         645 => x"6ff09ffb",
         646 => x"3357f600",
         647 => x"b396b600",
         648 => x"b366d700",
         649 => x"3357fe00",
         650 => x"331ebe00",
         651 => x"b357f300",
         652 => x"b3e7c701",
         653 => x"13de0601",
         654 => x"335fc703",
         655 => x"13980601",
         656 => x"13580801",
         657 => x"3316b600",
         658 => x"3377c703",
         659 => x"b30ee803",
         660 => x"13150701",
         661 => x"13d70701",
         662 => x"3367a700",
         663 => x"13050f00",
         664 => x"637ed701",
         665 => x"3387e600",
         666 => x"1305ffff",
         667 => x"6368d700",
         668 => x"6376d701",
         669 => x"1305efff",
         670 => x"3307d700",
         671 => x"3307d741",
         672 => x"b35ec703",
         673 => x"93970701",
         674 => x"93d70701",
         675 => x"3377c703",
         676 => x"3308d803",
         677 => x"13170701",
         678 => x"b3e7e700",
         679 => x"13870e00",
         680 => x"63fe0701",
         681 => x"b387f600",
         682 => x"1387feff",
         683 => x"63e8d700",
         684 => x"63f60701",
         685 => x"1387eeff",
         686 => x"b387d700",
         687 => x"13150501",
         688 => x"b70e0100",
         689 => x"3365e500",
         690 => x"9386feff",
         691 => x"3377d500",
         692 => x"b3870741",
         693 => x"b376d600",
         694 => x"13580501",
         695 => x"13560601",
         696 => x"330ed702",
         697 => x"b306d802",
         698 => x"3307c702",
         699 => x"3308c802",
         700 => x"3306d700",
         701 => x"13570e01",
         702 => x"3307c700",
         703 => x"6374d700",
         704 => x"3308d801",
         705 => x"93560701",
         706 => x"b3860601",
         707 => x"63e6d702",
         708 => x"e394d7ce",
         709 => x"b7070100",
         710 => x"9387f7ff",
         711 => x"3377f700",
         712 => x"13170701",
         713 => x"337efe00",
         714 => x"3313b300",
         715 => x"3307c701",
         716 => x"93050000",
         717 => x"e374e3da",
         718 => x"1305f5ff",
         719 => x"6ff0dfcb",
         720 => x"93050000",
         721 => x"13050000",
         722 => x"6ff05fd9",
         723 => x"93080500",
         724 => x"13830500",
         725 => x"13070600",
         726 => x"13080500",
         727 => x"93870500",
         728 => x"63920628",
         729 => x"b7450000",
         730 => x"93858593",
         731 => x"6376c30e",
         732 => x"b7060100",
         733 => x"6378d60c",
         734 => x"93360610",
         735 => x"93b61600",
         736 => x"93963600",
         737 => x"3355d600",
         738 => x"b385a500",
         739 => x"83c50500",
         740 => x"13050002",
         741 => x"b386d500",
         742 => x"b305d540",
         743 => x"630cd500",
         744 => x"b317b300",
         745 => x"b3d6d800",
         746 => x"3317b600",
         747 => x"b3e7f600",
         748 => x"3398b800",
         749 => x"93550701",
         750 => x"33d3b702",
         751 => x"13160701",
         752 => x"13560601",
         753 => x"b3f7b702",
         754 => x"13050300",
         755 => x"b3086602",
         756 => x"93960701",
         757 => x"93570801",
         758 => x"b3e7d700",
         759 => x"63fe1701",
         760 => x"b307f700",
         761 => x"1305f3ff",
         762 => x"63e8e700",
         763 => x"63f61701",
         764 => x"1305e3ff",
         765 => x"b387e700",
         766 => x"b3871741",
         767 => x"b3d8b702",
         768 => x"13180801",
         769 => x"13580801",
         770 => x"b3f7b702",
         771 => x"b3061603",
         772 => x"93970701",
         773 => x"3368f800",
         774 => x"93870800",
         775 => x"637cd800",
         776 => x"33080701",
         777 => x"9387f8ff",
         778 => x"6366e800",
         779 => x"6374d800",
         780 => x"9387e8ff",
         781 => x"13150501",
         782 => x"3365f500",
         783 => x"93050000",
         784 => x"67800000",
         785 => x"37050001",
         786 => x"93068001",
         787 => x"e37ca6f2",
         788 => x"93060001",
         789 => x"6ff01ff3",
         790 => x"93060000",
         791 => x"630c0600",
         792 => x"b7070100",
         793 => x"6370f60c",
         794 => x"93360610",
         795 => x"93b61600",
         796 => x"93963600",
         797 => x"b357d600",
         798 => x"b385f500",
         799 => x"83c70500",
         800 => x"b387d700",
         801 => x"93060002",
         802 => x"b385f640",
         803 => x"6396f60a",
         804 => x"b307c340",
         805 => x"93051000",
         806 => x"93580701",
         807 => x"33de1703",
         808 => x"13160701",
         809 => x"13560601",
         810 => x"93560801",
         811 => x"b3f71703",
         812 => x"13050e00",
         813 => x"3303c603",
         814 => x"93970701",
         815 => x"b3e7f600",
         816 => x"63fe6700",
         817 => x"b307f700",
         818 => x"1305feff",
         819 => x"63e8e700",
         820 => x"63f66700",
         821 => x"1305eeff",
         822 => x"b387e700",
         823 => x"b3876740",
         824 => x"33d31703",
         825 => x"13180801",
         826 => x"13580801",
         827 => x"b3f71703",
         828 => x"b3066602",
         829 => x"93970701",
         830 => x"3368f800",
         831 => x"93070300",
         832 => x"637cd800",
         833 => x"33080701",
         834 => x"9307f3ff",
         835 => x"6366e800",
         836 => x"6374d800",
         837 => x"9307e3ff",
         838 => x"13150501",
         839 => x"3365f500",
         840 => x"67800000",
         841 => x"b7070001",
         842 => x"93068001",
         843 => x"e374f6f4",
         844 => x"93060001",
         845 => x"6ff01ff4",
         846 => x"3317b600",
         847 => x"b356f300",
         848 => x"13550701",
         849 => x"3313b300",
         850 => x"b3d7f800",
         851 => x"b3e76700",
         852 => x"33d3a602",
         853 => x"13160701",
         854 => x"13560601",
         855 => x"3398b800",
         856 => x"b3f6a602",
         857 => x"b3086602",
         858 => x"93950601",
         859 => x"93d60701",
         860 => x"b3e6b600",
         861 => x"93050300",
         862 => x"63fe1601",
         863 => x"b306d700",
         864 => x"9305f3ff",
         865 => x"63e8e600",
         866 => x"63f61601",
         867 => x"9305e3ff",
         868 => x"b386e600",
         869 => x"b3861641",
         870 => x"b3d8a602",
         871 => x"93970701",
         872 => x"93d70701",
         873 => x"b3f6a602",
         874 => x"33061603",
         875 => x"93960601",
         876 => x"b3e7d700",
         877 => x"93860800",
         878 => x"63fec700",
         879 => x"b307f700",
         880 => x"9386f8ff",
         881 => x"63e8e700",
         882 => x"63f6c700",
         883 => x"9386e8ff",
         884 => x"b387e700",
         885 => x"93950501",
         886 => x"b387c740",
         887 => x"b3e5d500",
         888 => x"6ff09feb",
         889 => x"63e6d518",
         890 => x"b7070100",
         891 => x"63f4f604",
         892 => x"13b70610",
         893 => x"13371700",
         894 => x"13173700",
         895 => x"b7470000",
         896 => x"b3d5e600",
         897 => x"93878793",
         898 => x"b387b700",
         899 => x"83c70700",
         900 => x"b387e700",
         901 => x"13070002",
         902 => x"b305f740",
         903 => x"6316f702",
         904 => x"13051000",
         905 => x"e3ee66e0",
         906 => x"33b5c800",
         907 => x"13351500",
         908 => x"67800000",
         909 => x"b7070001",
         910 => x"13078001",
         911 => x"e3f0f6fc",
         912 => x"13070001",
         913 => x"6ff09ffb",
         914 => x"3357f600",
         915 => x"b396b600",
         916 => x"b366d700",
         917 => x"3357f300",
         918 => x"3313b300",
         919 => x"b3d7f800",
         920 => x"b3e76700",
         921 => x"13d30601",
         922 => x"b35e6702",
         923 => x"13980601",
         924 => x"13580801",
         925 => x"3316b600",
         926 => x"33776702",
         927 => x"330ed803",
         928 => x"13150701",
         929 => x"13d70701",
         930 => x"3367a700",
         931 => x"13850e00",
         932 => x"637ec701",
         933 => x"3387e600",
         934 => x"1385feff",
         935 => x"6368d700",
         936 => x"6376c701",
         937 => x"1385eeff",
         938 => x"3307d700",
         939 => x"3307c741",
         940 => x"335e6702",
         941 => x"93970701",
         942 => x"93d70701",
         943 => x"33776702",
         944 => x"3308c803",
         945 => x"13170701",
         946 => x"b3e7e700",
         947 => x"13070e00",
         948 => x"63fe0701",
         949 => x"b387f600",
         950 => x"1307feff",
         951 => x"63e8d700",
         952 => x"63f60701",
         953 => x"1307eeff",
         954 => x"b387d700",
         955 => x"13150501",
         956 => x"370e0100",
         957 => x"3365e500",
         958 => x"9306feff",
         959 => x"3377d500",
         960 => x"b3870741",
         961 => x"b376d600",
         962 => x"13580501",
         963 => x"13560601",
         964 => x"3303d702",
         965 => x"b306d802",
         966 => x"3307c702",
         967 => x"3308c802",
         968 => x"3306d700",
         969 => x"13570301",
         970 => x"3307c700",
         971 => x"6374d700",
         972 => x"3308c801",
         973 => x"93560701",
         974 => x"b3860601",
         975 => x"63e6d702",
         976 => x"e39ed7ce",
         977 => x"b7070100",
         978 => x"9387f7ff",
         979 => x"3377f700",
         980 => x"13170701",
         981 => x"3373f300",
         982 => x"b398b800",
         983 => x"33076700",
         984 => x"93050000",
         985 => x"e3fee8cc",
         986 => x"1305f5ff",
         987 => x"6ff01fcd",
         988 => x"93050000",
         989 => x"13050000",
         990 => x"67800000",
         991 => x"13080600",
         992 => x"93070500",
         993 => x"13870500",
         994 => x"63960620",
         995 => x"b7480000",
         996 => x"93888893",
         997 => x"63fcc50c",
         998 => x"b7060100",
         999 => x"637ed60a",
        1000 => x"93360610",
        1001 => x"93b61600",
        1002 => x"93963600",
        1003 => x"3353d600",
        1004 => x"b3886800",
        1005 => x"83c80800",
        1006 => x"13030002",
        1007 => x"b386d800",
        1008 => x"b308d340",
        1009 => x"630cd300",
        1010 => x"33971501",
        1011 => x"b356d500",
        1012 => x"33181601",
        1013 => x"33e7e600",
        1014 => x"b3171501",
        1015 => x"13560801",
        1016 => x"b356c702",
        1017 => x"13150801",
        1018 => x"13550501",
        1019 => x"3377c702",
        1020 => x"b386a602",
        1021 => x"93150701",
        1022 => x"13d70701",
        1023 => x"3367b700",
        1024 => x"637ad700",
        1025 => x"3307e800",
        1026 => x"63660701",
        1027 => x"6374d700",
        1028 => x"33070701",
        1029 => x"3307d740",
        1030 => x"b356c702",
        1031 => x"3377c702",
        1032 => x"b386a602",
        1033 => x"93970701",
        1034 => x"13170701",
        1035 => x"93d70701",
        1036 => x"b3e7e700",
        1037 => x"63fad700",
        1038 => x"b307f800",
        1039 => x"63e60701",
        1040 => x"63f4d700",
        1041 => x"b3870701",
        1042 => x"b387d740",
        1043 => x"33d51701",
        1044 => x"93050000",
        1045 => x"67800000",
        1046 => x"37030001",
        1047 => x"93068001",
        1048 => x"e37666f4",
        1049 => x"93060001",
        1050 => x"6ff05ff4",
        1051 => x"93060000",
        1052 => x"630c0600",
        1053 => x"37070100",
        1054 => x"637ee606",
        1055 => x"93360610",
        1056 => x"93b61600",
        1057 => x"93963600",
        1058 => x"3357d600",
        1059 => x"b388e800",
        1060 => x"03c70800",
        1061 => x"3307d700",
        1062 => x"93060002",
        1063 => x"b388e640",
        1064 => x"6394e606",
        1065 => x"3387c540",
        1066 => x"93550801",
        1067 => x"3356b702",
        1068 => x"13150801",
        1069 => x"13550501",
        1070 => x"93d60701",
        1071 => x"3377b702",
        1072 => x"3306a602",
        1073 => x"13170701",
        1074 => x"33e7e600",
        1075 => x"637ac700",
        1076 => x"3307e800",
        1077 => x"63660701",
        1078 => x"6374c700",
        1079 => x"33070701",
        1080 => x"3307c740",
        1081 => x"b356b702",
        1082 => x"3377b702",
        1083 => x"b386a602",
        1084 => x"6ff05ff3",
        1085 => x"37070001",
        1086 => x"93068001",
        1087 => x"e376e6f8",
        1088 => x"93060001",
        1089 => x"6ff05ff8",
        1090 => x"33181601",
        1091 => x"b3d6e500",
        1092 => x"b3171501",
        1093 => x"b3951501",
        1094 => x"3357e500",
        1095 => x"13550801",
        1096 => x"3367b700",
        1097 => x"b3d5a602",
        1098 => x"13130801",
        1099 => x"13530301",
        1100 => x"b3f6a602",
        1101 => x"b3856502",
        1102 => x"13960601",
        1103 => x"93560701",
        1104 => x"b3e6c600",
        1105 => x"63fab600",
        1106 => x"b306d800",
        1107 => x"63e60601",
        1108 => x"63f4b600",
        1109 => x"b3860601",
        1110 => x"b386b640",
        1111 => x"33d6a602",
        1112 => x"13170701",
        1113 => x"13570701",
        1114 => x"b3f6a602",
        1115 => x"33066602",
        1116 => x"93960601",
        1117 => x"3367d700",
        1118 => x"637ac700",
        1119 => x"3307e800",
        1120 => x"63660701",
        1121 => x"6374c700",
        1122 => x"33070701",
        1123 => x"3307c740",
        1124 => x"6ff09ff1",
        1125 => x"63e4d51c",
        1126 => x"37080100",
        1127 => x"63fe0605",
        1128 => x"13b80610",
        1129 => x"13381800",
        1130 => x"13183800",
        1131 => x"b7480000",
        1132 => x"33d30601",
        1133 => x"93888893",
        1134 => x"b3886800",
        1135 => x"83c80800",
        1136 => x"13030002",
        1137 => x"b3880801",
        1138 => x"33081341",
        1139 => x"63101305",
        1140 => x"63e4b600",
        1141 => x"636cc500",
        1142 => x"3306c540",
        1143 => x"b386d540",
        1144 => x"3337c500",
        1145 => x"93070600",
        1146 => x"3387e640",
        1147 => x"13850700",
        1148 => x"93050700",
        1149 => x"67800000",
        1150 => x"b7080001",
        1151 => x"13088001",
        1152 => x"e3f616fb",
        1153 => x"13080001",
        1154 => x"6ff05ffa",
        1155 => x"b3571601",
        1156 => x"b3960601",
        1157 => x"b3e6d700",
        1158 => x"33d71501",
        1159 => x"13de0601",
        1160 => x"335fc703",
        1161 => x"13930601",
        1162 => x"13530301",
        1163 => x"b3970501",
        1164 => x"b3551501",
        1165 => x"b3e5f500",
        1166 => x"93d70501",
        1167 => x"33160601",
        1168 => x"33150501",
        1169 => x"3377c703",
        1170 => x"b30ee303",
        1171 => x"13170701",
        1172 => x"b3e7e700",
        1173 => x"13070f00",
        1174 => x"63fed701",
        1175 => x"b387f600",
        1176 => x"1307ffff",
        1177 => x"63e8d700",
        1178 => x"63f6d701",
        1179 => x"1307efff",
        1180 => x"b387d700",
        1181 => x"b387d741",
        1182 => x"b3dec703",
        1183 => x"93950501",
        1184 => x"93d50501",
        1185 => x"b3f7c703",
        1186 => x"138e0e00",
        1187 => x"3303d303",
        1188 => x"93970701",
        1189 => x"b3e5f500",
        1190 => x"63fe6500",
        1191 => x"b385b600",
        1192 => x"138efeff",
        1193 => x"63e8d500",
        1194 => x"63f66500",
        1195 => x"138eeeff",
        1196 => x"b385d500",
        1197 => x"93170701",
        1198 => x"370f0100",
        1199 => x"b3e7c701",
        1200 => x"b3856540",
        1201 => x"1303ffff",
        1202 => x"33f76700",
        1203 => x"135e0601",
        1204 => x"93d70701",
        1205 => x"33736600",
        1206 => x"b30e6702",
        1207 => x"33836702",
        1208 => x"3307c703",
        1209 => x"b387c703",
        1210 => x"330e6700",
        1211 => x"13d70e01",
        1212 => x"3307c701",
        1213 => x"63746700",
        1214 => x"b387e701",
        1215 => x"13530701",
        1216 => x"b307f300",
        1217 => x"37030100",
        1218 => x"1303f3ff",
        1219 => x"33776700",
        1220 => x"13170701",
        1221 => x"b3fe6e00",
        1222 => x"3307d701",
        1223 => x"63e6f500",
        1224 => x"639ef500",
        1225 => x"637ce500",
        1226 => x"3306c740",
        1227 => x"3333c700",
        1228 => x"b306d300",
        1229 => x"13070600",
        1230 => x"b387d740",
        1231 => x"3307e540",
        1232 => x"3335e500",
        1233 => x"b385f540",
        1234 => x"b385a540",
        1235 => x"b3981501",
        1236 => x"33570701",
        1237 => x"33e5e800",
        1238 => x"b3d50501",
        1239 => x"67800000",
        1240 => x"13030500",
        1241 => x"630a0600",
        1242 => x"2300b300",
        1243 => x"1306f6ff",
        1244 => x"13031300",
        1245 => x"e31a06fe",
        1246 => x"67800000",
        1247 => x"13030500",
        1248 => x"630e0600",
        1249 => x"83830500",
        1250 => x"23007300",
        1251 => x"1306f6ff",
        1252 => x"13031300",
        1253 => x"93851500",
        1254 => x"e31606fe",
        1255 => x"67800000",
        1256 => x"630c0602",
        1257 => x"13030500",
        1258 => x"93061000",
        1259 => x"636ab500",
        1260 => x"9306f0ff",
        1261 => x"1307f6ff",
        1262 => x"3303e300",
        1263 => x"b385e500",
        1264 => x"83830500",
        1265 => x"23007300",
        1266 => x"1306f6ff",
        1267 => x"3303d300",
        1268 => x"b385d500",
        1269 => x"e31606fe",
        1270 => x"67800000",
        1271 => x"6f000000",
        1272 => x"130101ff",
        1273 => x"23248100",
        1274 => x"13040000",
        1275 => x"23229100",
        1276 => x"23202101",
        1277 => x"23261100",
        1278 => x"93040500",
        1279 => x"13090400",
        1280 => x"93070400",
        1281 => x"732410c8",
        1282 => x"732910c0",
        1283 => x"f32710c8",
        1284 => x"e31af4fe",
        1285 => x"37460f00",
        1286 => x"13060624",
        1287 => x"93060000",
        1288 => x"13050900",
        1289 => x"93050400",
        1290 => x"eff05fb5",
        1291 => x"37460f00",
        1292 => x"23a4a400",
        1293 => x"93050400",
        1294 => x"13050900",
        1295 => x"13060624",
        1296 => x"93060000",
        1297 => x"eff08ff0",
        1298 => x"8320c100",
        1299 => x"03248100",
        1300 => x"23a0a400",
        1301 => x"23a2b400",
        1302 => x"03290100",
        1303 => x"83244100",
        1304 => x"13050000",
        1305 => x"13010101",
        1306 => x"67800000",
        1307 => x"13050000",
        1308 => x"67800000",
        1309 => x"13050000",
        1310 => x"67800000",
        1311 => x"130101ff",
        1312 => x"23202101",
        1313 => x"23261100",
        1314 => x"13090600",
        1315 => x"6356c002",
        1316 => x"23248100",
        1317 => x"23229100",
        1318 => x"13840500",
        1319 => x"b384c500",
        1320 => x"03450400",
        1321 => x"13041400",
        1322 => x"efe05fbd",
        1323 => x"e39a84fe",
        1324 => x"03248100",
        1325 => x"83244100",
        1326 => x"8320c100",
        1327 => x"13050900",
        1328 => x"03290100",
        1329 => x"13010101",
        1330 => x"67800000",
        1331 => x"130101ff",
        1332 => x"23202101",
        1333 => x"23261100",
        1334 => x"13090600",
        1335 => x"6356c002",
        1336 => x"23248100",
        1337 => x"23229100",
        1338 => x"13840500",
        1339 => x"b384c500",
        1340 => x"efe09fb8",
        1341 => x"13041400",
        1342 => x"a30fa4fe",
        1343 => x"e39a84fe",
        1344 => x"03248100",
        1345 => x"83244100",
        1346 => x"8320c100",
        1347 => x"13050900",
        1348 => x"03290100",
        1349 => x"13010101",
        1350 => x"67800000",
        1351 => x"13051000",
        1352 => x"67800000",
        1353 => x"130101ff",
        1354 => x"23261100",
        1355 => x"ef00d060",
        1356 => x"8320c100",
        1357 => x"93076001",
        1358 => x"2320f500",
        1359 => x"1305f0ff",
        1360 => x"13010101",
        1361 => x"67800000",
        1362 => x"1305f0ff",
        1363 => x"67800000",
        1364 => x"b7270000",
        1365 => x"23a2f500",
        1366 => x"13050000",
        1367 => x"67800000",
        1368 => x"13051000",
        1369 => x"67800000",
        1370 => x"13050000",
        1371 => x"67800000",
        1372 => x"130101fe",
        1373 => x"2324c100",
        1374 => x"2326d100",
        1375 => x"2328e100",
        1376 => x"232af100",
        1377 => x"232c0101",
        1378 => x"232e1101",
        1379 => x"1305f0ff",
        1380 => x"13010102",
        1381 => x"67800000",
        1382 => x"130101ff",
        1383 => x"23261100",
        1384 => x"ef009059",
        1385 => x"8320c100",
        1386 => x"9307a000",
        1387 => x"2320f500",
        1388 => x"1305f0ff",
        1389 => x"13010101",
        1390 => x"67800000",
        1391 => x"130101ff",
        1392 => x"23261100",
        1393 => x"ef005057",
        1394 => x"8320c100",
        1395 => x"93072000",
        1396 => x"2320f500",
        1397 => x"1305f0ff",
        1398 => x"13010101",
        1399 => x"67800000",
        1400 => x"b7270000",
        1401 => x"23a2f500",
        1402 => x"13050000",
        1403 => x"67800000",
        1404 => x"130101ff",
        1405 => x"23261100",
        1406 => x"ef001054",
        1407 => x"8320c100",
        1408 => x"9307f001",
        1409 => x"2320f500",
        1410 => x"1305f0ff",
        1411 => x"13010101",
        1412 => x"67800000",
        1413 => x"130101ff",
        1414 => x"23261100",
        1415 => x"ef00d051",
        1416 => x"8320c100",
        1417 => x"9307b000",
        1418 => x"2320f500",
        1419 => x"1305f0ff",
        1420 => x"13010101",
        1421 => x"67800000",
        1422 => x"130101ff",
        1423 => x"23261100",
        1424 => x"ef00904f",
        1425 => x"8320c100",
        1426 => x"9307c000",
        1427 => x"2320f500",
        1428 => x"1305f0ff",
        1429 => x"13010101",
        1430 => x"67800000",
        1431 => x"03a7c187",
        1432 => x"b7870020",
        1433 => x"93870700",
        1434 => x"93060040",
        1435 => x"b387d740",
        1436 => x"630c0700",
        1437 => x"3305a700",
        1438 => x"63e2a702",
        1439 => x"23aea186",
        1440 => x"13050700",
        1441 => x"67800000",
        1442 => x"9386819c",
        1443 => x"1387819c",
        1444 => x"23aed186",
        1445 => x"3305a700",
        1446 => x"e3f2a7fe",
        1447 => x"130101ff",
        1448 => x"23261100",
        1449 => x"ef005049",
        1450 => x"8320c100",
        1451 => x"9307c000",
        1452 => x"2320f500",
        1453 => x"1307f0ff",
        1454 => x"13050700",
        1455 => x"13010101",
        1456 => x"67800000",
        1457 => x"370700f0",
        1458 => x"13070702",
        1459 => x"83274700",
        1460 => x"93f74700",
        1461 => x"e38c07fe",
        1462 => x"03258700",
        1463 => x"1375f50f",
        1464 => x"67800000",
        1465 => x"f32710fc",
        1466 => x"63960700",
        1467 => x"b7f7fa02",
        1468 => x"93870708",
        1469 => x"63060500",
        1470 => x"33d5a702",
        1471 => x"1305f5ff",
        1472 => x"b70700f0",
        1473 => x"23a6a702",
        1474 => x"23a0b702",
        1475 => x"67800000",
        1476 => x"370700f0",
        1477 => x"1375f50f",
        1478 => x"13070702",
        1479 => x"2324a700",
        1480 => x"83274700",
        1481 => x"93f70701",
        1482 => x"e38c07fe",
        1483 => x"67800000",
        1484 => x"630e0502",
        1485 => x"130101ff",
        1486 => x"23248100",
        1487 => x"23261100",
        1488 => x"13040500",
        1489 => x"03450500",
        1490 => x"630a0500",
        1491 => x"13041400",
        1492 => x"eff01ffc",
        1493 => x"03450400",
        1494 => x"e31a05fe",
        1495 => x"8320c100",
        1496 => x"03248100",
        1497 => x"13010101",
        1498 => x"67800000",
        1499 => x"67800000",
        1500 => x"130101f9",
        1501 => x"23229106",
        1502 => x"23202107",
        1503 => x"23261106",
        1504 => x"23248106",
        1505 => x"232e3105",
        1506 => x"232c4105",
        1507 => x"232a5105",
        1508 => x"23286105",
        1509 => x"23267105",
        1510 => x"23248105",
        1511 => x"23229105",
        1512 => x"2320a105",
        1513 => x"13090500",
        1514 => x"93840500",
        1515 => x"232c0100",
        1516 => x"232e0100",
        1517 => x"23200102",
        1518 => x"23220102",
        1519 => x"23240102",
        1520 => x"23260102",
        1521 => x"23280102",
        1522 => x"232a0102",
        1523 => x"232c0102",
        1524 => x"232e0102",
        1525 => x"732410fc",
        1526 => x"63160400",
        1527 => x"37f4fa02",
        1528 => x"13040408",
        1529 => x"97f2ffff",
        1530 => x"938242b0",
        1531 => x"73905230",
        1532 => x"37c50100",
        1533 => x"93050004",
        1534 => x"13050520",
        1535 => x"eff09fee",
        1536 => x"b7270000",
        1537 => x"93870771",
        1538 => x"b356f402",
        1539 => x"13561400",
        1540 => x"370700f0",
        1541 => x"1306f6ff",
        1542 => x"b7170300",
        1543 => x"2326c708",
        1544 => x"130e1001",
        1545 => x"938707d4",
        1546 => x"2320c709",
        1547 => x"370600f0",
        1548 => x"37230000",
        1549 => x"1303f370",
        1550 => x"37581200",
        1551 => x"130808f8",
        1552 => x"b70800f0",
        1553 => x"370500f0",
        1554 => x"b70500f0",
        1555 => x"3357f402",
        1556 => x"9387f6ff",
        1557 => x"2328f60a",
        1558 => x"2326660a",
        1559 => x"2320c60b",
        1560 => x"93078070",
        1561 => x"23a0f806",
        1562 => x"b3570403",
        1563 => x"1307f7ff",
        1564 => x"13170701",
        1565 => x"13678700",
        1566 => x"2320e504",
        1567 => x"1307a007",
        1568 => x"9387f7ff",
        1569 => x"93970701",
        1570 => x"93e7c700",
        1571 => x"23a8f504",
        1572 => x"b70700f0",
        1573 => x"23ace700",
        1574 => x"93020008",
        1575 => x"73904230",
        1576 => x"b7220000",
        1577 => x"93828280",
        1578 => x"73900230",
        1579 => x"b7490000",
        1580 => x"138589a5",
        1581 => x"eff0dfe7",
        1582 => x"1304f9ff",
        1583 => x"63522003",
        1584 => x"1309f0ff",
        1585 => x"03a50400",
        1586 => x"1304f4ff",
        1587 => x"93844400",
        1588 => x"eff01fe6",
        1589 => x"138589a5",
        1590 => x"eff09fe5",
        1591 => x"e31424ff",
        1592 => x"37450000",
        1593 => x"1305c5a5",
        1594 => x"37f9eeee",
        1595 => x"b7faeeee",
        1596 => x"b7090010",
        1597 => x"37140000",
        1598 => x"eff09fe3",
        1599 => x"374b0000",
        1600 => x"9389f9ff",
        1601 => x"1309f9ee",
        1602 => x"938aeaee",
        1603 => x"130404e1",
        1604 => x"93040000",
        1605 => x"b71b0000",
        1606 => x"938b0b2c",
        1607 => x"130af000",
        1608 => x"6f00c000",
        1609 => x"938bfbff",
        1610 => x"63840b18",
        1611 => x"93050000",
        1612 => x"13058100",
        1613 => x"ef00902a",
        1614 => x"e31605fe",
        1615 => x"032c8100",
        1616 => x"8325c100",
        1617 => x"13060400",
        1618 => x"9357cc01",
        1619 => x"13974500",
        1620 => x"b367f700",
        1621 => x"b3f73701",
        1622 => x"33773c01",
        1623 => x"13d5f541",
        1624 => x"13d88501",
        1625 => x"3307f700",
        1626 => x"33070701",
        1627 => x"9377d500",
        1628 => x"3307f700",
        1629 => x"33774703",
        1630 => x"937725ff",
        1631 => x"93860400",
        1632 => x"13050c00",
        1633 => x"938bfbff",
        1634 => x"3307f700",
        1635 => x"b307ec40",
        1636 => x"1357f741",
        1637 => x"3338fc00",
        1638 => x"3387e540",
        1639 => x"33070741",
        1640 => x"b3885703",
        1641 => x"33072703",
        1642 => x"33b82703",
        1643 => x"33071701",
        1644 => x"b3872703",
        1645 => x"33070701",
        1646 => x"1358f741",
        1647 => x"13783800",
        1648 => x"b307f800",
        1649 => x"33b80701",
        1650 => x"3307e800",
        1651 => x"1318e701",
        1652 => x"93d72700",
        1653 => x"b367f800",
        1654 => x"13582740",
        1655 => x"93184800",
        1656 => x"13d3c701",
        1657 => x"33e36800",
        1658 => x"33733301",
        1659 => x"b3f83701",
        1660 => x"135e8801",
        1661 => x"1357f741",
        1662 => x"b3886800",
        1663 => x"b388c801",
        1664 => x"1373d700",
        1665 => x"b3886800",
        1666 => x"b3f84803",
        1667 => x"137727ff",
        1668 => x"939c4700",
        1669 => x"b38cfc40",
        1670 => x"939c2c00",
        1671 => x"b30c9c41",
        1672 => x"b388e800",
        1673 => x"33871741",
        1674 => x"93d8f841",
        1675 => x"33b3e700",
        1676 => x"33081841",
        1677 => x"33086840",
        1678 => x"33082803",
        1679 => x"33035703",
        1680 => x"b3382703",
        1681 => x"33086800",
        1682 => x"33072703",
        1683 => x"33081801",
        1684 => x"9358f841",
        1685 => x"93f83800",
        1686 => x"3387e800",
        1687 => x"b3381701",
        1688 => x"b3880801",
        1689 => x"9398e801",
        1690 => x"13572700",
        1691 => x"33e7e800",
        1692 => x"13184700",
        1693 => x"3307e840",
        1694 => x"13172700",
        1695 => x"338de740",
        1696 => x"efe05fc5",
        1697 => x"83260101",
        1698 => x"13070500",
        1699 => x"13880c00",
        1700 => x"93070d00",
        1701 => x"13060c00",
        1702 => x"9305cba8",
        1703 => x"13058101",
        1704 => x"ef00c045",
        1705 => x"13058101",
        1706 => x"eff09fc8",
        1707 => x"e3900be8",
        1708 => x"73001000",
        1709 => x"b70700f0",
        1710 => x"9306f00f",
        1711 => x"23a4d706",
        1712 => x"370700f0",
        1713 => x"83260704",
        1714 => x"13060009",
        1715 => x"b70700f0",
        1716 => x"93e60630",
        1717 => x"2320d704",
        1718 => x"2324c704",
        1719 => x"83a60705",
        1720 => x"13e70630",
        1721 => x"23a8e704",
        1722 => x"23acc704",
        1723 => x"6ff09fe2",
        1724 => x"130101ff",
        1725 => x"23248100",
        1726 => x"23261100",
        1727 => x"93070000",
        1728 => x"13040500",
        1729 => x"63880700",
        1730 => x"93050000",
        1731 => x"97000000",
        1732 => x"e7000000",
        1733 => x"83a70188",
        1734 => x"63840700",
        1735 => x"e7800700",
        1736 => x"13050400",
        1737 => x"eff09f8b",
        1738 => x"13050000",
        1739 => x"67800000",
        1740 => x"130101ff",
        1741 => x"23248100",
        1742 => x"23261100",
        1743 => x"13040500",
        1744 => x"2316b500",
        1745 => x"2317c500",
        1746 => x"23200500",
        1747 => x"23220500",
        1748 => x"23240500",
        1749 => x"23220506",
        1750 => x"23280500",
        1751 => x"232a0500",
        1752 => x"232c0500",
        1753 => x"13068000",
        1754 => x"93050000",
        1755 => x"1305c505",
        1756 => x"eff00fff",
        1757 => x"b7270000",
        1758 => x"9387c7f6",
        1759 => x"2322f402",
        1760 => x"b7270000",
        1761 => x"938747fc",
        1762 => x"2324f402",
        1763 => x"b7270000",
        1764 => x"93878704",
        1765 => x"2326f402",
        1766 => x"b7270000",
        1767 => x"9387070a",
        1768 => x"8320c100",
        1769 => x"23208402",
        1770 => x"2328f402",
        1771 => x"03248100",
        1772 => x"13010101",
        1773 => x"67800000",
        1774 => x"b7350000",
        1775 => x"37050020",
        1776 => x"13868181",
        1777 => x"93858551",
        1778 => x"13054502",
        1779 => x"6f00c021",
        1780 => x"83254500",
        1781 => x"130101ff",
        1782 => x"b7070020",
        1783 => x"23248100",
        1784 => x"23261100",
        1785 => x"93870709",
        1786 => x"13040500",
        1787 => x"6384f500",
        1788 => x"ef109012",
        1789 => x"83258400",
        1790 => x"9387818f",
        1791 => x"6386f500",
        1792 => x"13050400",
        1793 => x"ef105011",
        1794 => x"8325c400",
        1795 => x"93870196",
        1796 => x"638cf500",
        1797 => x"13050400",
        1798 => x"03248100",
        1799 => x"8320c100",
        1800 => x"13010101",
        1801 => x"6f10500f",
        1802 => x"8320c100",
        1803 => x"03248100",
        1804 => x"13010101",
        1805 => x"67800000",
        1806 => x"b7270000",
        1807 => x"37050020",
        1808 => x"130101ff",
        1809 => x"938787bb",
        1810 => x"13060000",
        1811 => x"93054000",
        1812 => x"13050509",
        1813 => x"23261100",
        1814 => x"23a0f188",
        1815 => x"eff05fed",
        1816 => x"13061000",
        1817 => x"93059000",
        1818 => x"1385818f",
        1819 => x"eff05fec",
        1820 => x"8320c100",
        1821 => x"13062000",
        1822 => x"93052001",
        1823 => x"13850196",
        1824 => x"13010101",
        1825 => x"6ff0dfea",
        1826 => x"13050000",
        1827 => x"67800000",
        1828 => x"83a70188",
        1829 => x"130101ff",
        1830 => x"23202101",
        1831 => x"23261100",
        1832 => x"23248100",
        1833 => x"23229100",
        1834 => x"13090500",
        1835 => x"63940700",
        1836 => x"eff09ff8",
        1837 => x"93848181",
        1838 => x"03a48400",
        1839 => x"83a74400",
        1840 => x"9387f7ff",
        1841 => x"63d80702",
        1842 => x"83a70400",
        1843 => x"6390070c",
        1844 => x"9305c01a",
        1845 => x"13050900",
        1846 => x"ef001009",
        1847 => x"13040500",
        1848 => x"63140508",
        1849 => x"23a00400",
        1850 => x"9307c000",
        1851 => x"2320f900",
        1852 => x"6f004005",
        1853 => x"0317c400",
        1854 => x"63140706",
        1855 => x"b707ffff",
        1856 => x"93871700",
        1857 => x"23220406",
        1858 => x"23200400",
        1859 => x"23220400",
        1860 => x"23240400",
        1861 => x"2326f400",
        1862 => x"23280400",
        1863 => x"232a0400",
        1864 => x"232c0400",
        1865 => x"13068000",
        1866 => x"93050000",
        1867 => x"1305c405",
        1868 => x"eff00fe3",
        1869 => x"232a0402",
        1870 => x"232c0402",
        1871 => x"23240404",
        1872 => x"23260404",
        1873 => x"8320c100",
        1874 => x"13050400",
        1875 => x"03248100",
        1876 => x"83244100",
        1877 => x"03290100",
        1878 => x"13010101",
        1879 => x"67800000",
        1880 => x"13048406",
        1881 => x"6ff0dff5",
        1882 => x"93074000",
        1883 => x"23200500",
        1884 => x"2322f500",
        1885 => x"1305c500",
        1886 => x"2324a400",
        1887 => x"1306001a",
        1888 => x"93050000",
        1889 => x"eff0cfdd",
        1890 => x"23a08400",
        1891 => x"83a40400",
        1892 => x"6ff09ff2",
        1893 => x"83270502",
        1894 => x"639e0700",
        1895 => x"b7270000",
        1896 => x"938707bd",
        1897 => x"2320f502",
        1898 => x"83a70188",
        1899 => x"63940700",
        1900 => x"6ff09fe8",
        1901 => x"67800000",
        1902 => x"67800000",
        1903 => x"67800000",
        1904 => x"b7250000",
        1905 => x"13868181",
        1906 => x"938585b2",
        1907 => x"13050000",
        1908 => x"6f008001",
        1909 => x"b7250000",
        1910 => x"13868181",
        1911 => x"938585c8",
        1912 => x"13050000",
        1913 => x"6f004000",
        1914 => x"130101fd",
        1915 => x"23248102",
        1916 => x"23202103",
        1917 => x"232e3101",
        1918 => x"232c4101",
        1919 => x"23286101",
        1920 => x"23267101",
        1921 => x"23261102",
        1922 => x"23229102",
        1923 => x"232a5101",
        1924 => x"93090500",
        1925 => x"138a0500",
        1926 => x"13040600",
        1927 => x"13090000",
        1928 => x"130b1000",
        1929 => x"930bf0ff",
        1930 => x"83248400",
        1931 => x"832a4400",
        1932 => x"938afaff",
        1933 => x"63de0a02",
        1934 => x"03240400",
        1935 => x"e31604fe",
        1936 => x"8320c102",
        1937 => x"03248102",
        1938 => x"83244102",
        1939 => x"8329c101",
        1940 => x"032a8101",
        1941 => x"832a4101",
        1942 => x"032b0101",
        1943 => x"832bc100",
        1944 => x"13050900",
        1945 => x"03290102",
        1946 => x"13010103",
        1947 => x"67800000",
        1948 => x"83d7c400",
        1949 => x"637efb00",
        1950 => x"8397e400",
        1951 => x"638a7701",
        1952 => x"93850400",
        1953 => x"13850900",
        1954 => x"e7000a00",
        1955 => x"3369a900",
        1956 => x"93848406",
        1957 => x"6ff0dff9",
        1958 => x"130101f6",
        1959 => x"232af108",
        1960 => x"b7070080",
        1961 => x"9387f7ff",
        1962 => x"232ef100",
        1963 => x"2328f100",
        1964 => x"b707ffff",
        1965 => x"2326d108",
        1966 => x"2324b100",
        1967 => x"232cb100",
        1968 => x"93878720",
        1969 => x"9306c108",
        1970 => x"93058100",
        1971 => x"232e1106",
        1972 => x"232af100",
        1973 => x"2328e108",
        1974 => x"232c0109",
        1975 => x"232e1109",
        1976 => x"2322d100",
        1977 => x"ef00d037",
        1978 => x"83278100",
        1979 => x"23800700",
        1980 => x"8320c107",
        1981 => x"1301010a",
        1982 => x"67800000",
        1983 => x"130101f6",
        1984 => x"232af108",
        1985 => x"b7070080",
        1986 => x"9387f7ff",
        1987 => x"232ef100",
        1988 => x"2328f100",
        1989 => x"b707ffff",
        1990 => x"93878720",
        1991 => x"232af100",
        1992 => x"2324a100",
        1993 => x"232ca100",
        1994 => x"03a54187",
        1995 => x"2324c108",
        1996 => x"2326d108",
        1997 => x"13860500",
        1998 => x"93068108",
        1999 => x"93058100",
        2000 => x"232e1106",
        2001 => x"2328e108",
        2002 => x"232c0109",
        2003 => x"232e1109",
        2004 => x"2322d100",
        2005 => x"ef00d030",
        2006 => x"83278100",
        2007 => x"23800700",
        2008 => x"8320c107",
        2009 => x"1301010a",
        2010 => x"67800000",
        2011 => x"130101ff",
        2012 => x"23248100",
        2013 => x"13840500",
        2014 => x"8395e500",
        2015 => x"23261100",
        2016 => x"ef008031",
        2017 => x"63400502",
        2018 => x"83274405",
        2019 => x"b387a700",
        2020 => x"232af404",
        2021 => x"8320c100",
        2022 => x"03248100",
        2023 => x"13010101",
        2024 => x"67800000",
        2025 => x"8357c400",
        2026 => x"37f7ffff",
        2027 => x"1307f7ff",
        2028 => x"b3f7e700",
        2029 => x"2316f400",
        2030 => x"6ff0dffd",
        2031 => x"13050000",
        2032 => x"67800000",
        2033 => x"83d7c500",
        2034 => x"130101fe",
        2035 => x"232c8100",
        2036 => x"232a9100",
        2037 => x"23282101",
        2038 => x"23263101",
        2039 => x"232e1100",
        2040 => x"93f70710",
        2041 => x"93040500",
        2042 => x"13840500",
        2043 => x"13090600",
        2044 => x"93890600",
        2045 => x"638a0700",
        2046 => x"8395e500",
        2047 => x"93062000",
        2048 => x"13060000",
        2049 => x"ef004024",
        2050 => x"8357c400",
        2051 => x"37f7ffff",
        2052 => x"1307f7ff",
        2053 => x"b3f7e700",
        2054 => x"8315e400",
        2055 => x"2316f400",
        2056 => x"03248101",
        2057 => x"8320c101",
        2058 => x"93860900",
        2059 => x"13060900",
        2060 => x"8329c100",
        2061 => x"03290101",
        2062 => x"13850400",
        2063 => x"83244101",
        2064 => x"13010102",
        2065 => x"6f00402a",
        2066 => x"130101ff",
        2067 => x"23248100",
        2068 => x"13840500",
        2069 => x"8395e500",
        2070 => x"23261100",
        2071 => x"ef00c01e",
        2072 => x"1307f0ff",
        2073 => x"8357c400",
        2074 => x"6312e502",
        2075 => x"37f7ffff",
        2076 => x"1307f7ff",
        2077 => x"b3f7e700",
        2078 => x"2316f400",
        2079 => x"8320c100",
        2080 => x"03248100",
        2081 => x"13010101",
        2082 => x"67800000",
        2083 => x"37170000",
        2084 => x"b3e7e700",
        2085 => x"2316f400",
        2086 => x"232aa404",
        2087 => x"6ff01ffe",
        2088 => x"8395e500",
        2089 => x"6f004000",
        2090 => x"130101ff",
        2091 => x"23248100",
        2092 => x"23229100",
        2093 => x"13040500",
        2094 => x"13850500",
        2095 => x"23261100",
        2096 => x"23a20188",
        2097 => x"eff04fc8",
        2098 => x"9307f0ff",
        2099 => x"6318f500",
        2100 => x"83a74188",
        2101 => x"63840700",
        2102 => x"2320f400",
        2103 => x"8320c100",
        2104 => x"03248100",
        2105 => x"83244100",
        2106 => x"13010101",
        2107 => x"67800000",
        2108 => x"83a74187",
        2109 => x"6388a714",
        2110 => x"8327c501",
        2111 => x"130101fe",
        2112 => x"232c8100",
        2113 => x"232e1100",
        2114 => x"232a9100",
        2115 => x"23282101",
        2116 => x"23263101",
        2117 => x"13040500",
        2118 => x"638a0704",
        2119 => x"83a7c700",
        2120 => x"638c0702",
        2121 => x"93040000",
        2122 => x"13090008",
        2123 => x"8327c401",
        2124 => x"83a7c700",
        2125 => x"b3879700",
        2126 => x"83a50700",
        2127 => x"639c050c",
        2128 => x"93844400",
        2129 => x"e39424ff",
        2130 => x"8327c401",
        2131 => x"13050400",
        2132 => x"83a5c700",
        2133 => x"ef008029",
        2134 => x"8327c401",
        2135 => x"83a50700",
        2136 => x"63860500",
        2137 => x"13050400",
        2138 => x"ef004028",
        2139 => x"83254401",
        2140 => x"63860500",
        2141 => x"13050400",
        2142 => x"ef004027",
        2143 => x"8325c401",
        2144 => x"63860500",
        2145 => x"13050400",
        2146 => x"ef004026",
        2147 => x"83250403",
        2148 => x"63860500",
        2149 => x"13050400",
        2150 => x"ef004025",
        2151 => x"83254403",
        2152 => x"63860500",
        2153 => x"13050400",
        2154 => x"ef004024",
        2155 => x"83258403",
        2156 => x"63860500",
        2157 => x"13050400",
        2158 => x"ef004023",
        2159 => x"83258404",
        2160 => x"63860500",
        2161 => x"13050400",
        2162 => x"ef004022",
        2163 => x"83254404",
        2164 => x"63860500",
        2165 => x"13050400",
        2166 => x"ef004021",
        2167 => x"8325c402",
        2168 => x"63860500",
        2169 => x"13050400",
        2170 => x"ef004020",
        2171 => x"83270402",
        2172 => x"638c0702",
        2173 => x"13050400",
        2174 => x"03248101",
        2175 => x"8320c101",
        2176 => x"83244101",
        2177 => x"03290101",
        2178 => x"8329c100",
        2179 => x"13010102",
        2180 => x"67800700",
        2181 => x"83a90500",
        2182 => x"13050400",
        2183 => x"ef00001d",
        2184 => x"93850900",
        2185 => x"6ff09ff1",
        2186 => x"8320c101",
        2187 => x"03248101",
        2188 => x"83244101",
        2189 => x"03290101",
        2190 => x"8329c100",
        2191 => x"13010102",
        2192 => x"67800000",
        2193 => x"67800000",
        2194 => x"130101ff",
        2195 => x"23248100",
        2196 => x"23229100",
        2197 => x"13040500",
        2198 => x"13850500",
        2199 => x"93050600",
        2200 => x"13860600",
        2201 => x"23261100",
        2202 => x"23a20188",
        2203 => x"eff0cfaf",
        2204 => x"9307f0ff",
        2205 => x"6318f500",
        2206 => x"83a74188",
        2207 => x"63840700",
        2208 => x"2320f400",
        2209 => x"8320c100",
        2210 => x"03248100",
        2211 => x"83244100",
        2212 => x"13010101",
        2213 => x"67800000",
        2214 => x"130101ff",
        2215 => x"23248100",
        2216 => x"23229100",
        2217 => x"13040500",
        2218 => x"13850500",
        2219 => x"93050600",
        2220 => x"13860600",
        2221 => x"23261100",
        2222 => x"23a20188",
        2223 => x"eff00fa1",
        2224 => x"9307f0ff",
        2225 => x"6318f500",
        2226 => x"83a74188",
        2227 => x"63840700",
        2228 => x"2320f400",
        2229 => x"8320c100",
        2230 => x"03248100",
        2231 => x"83244100",
        2232 => x"13010101",
        2233 => x"67800000",
        2234 => x"130101ff",
        2235 => x"23248100",
        2236 => x"23229100",
        2237 => x"13040500",
        2238 => x"13850500",
        2239 => x"93050600",
        2240 => x"13860600",
        2241 => x"23261100",
        2242 => x"23a20188",
        2243 => x"eff00f97",
        2244 => x"9307f0ff",
        2245 => x"6318f500",
        2246 => x"83a74188",
        2247 => x"63840700",
        2248 => x"2320f400",
        2249 => x"8320c100",
        2250 => x"03248100",
        2251 => x"83244100",
        2252 => x"13010101",
        2253 => x"67800000",
        2254 => x"03a54187",
        2255 => x"67800000",
        2256 => x"130101ff",
        2257 => x"23248100",
        2258 => x"23229100",
        2259 => x"37440000",
        2260 => x"b7440000",
        2261 => x"9387c4be",
        2262 => x"1304c4be",
        2263 => x"3304f440",
        2264 => x"23202101",
        2265 => x"23261100",
        2266 => x"13542440",
        2267 => x"9384c4be",
        2268 => x"13090000",
        2269 => x"63108904",
        2270 => x"b7440000",
        2271 => x"37440000",
        2272 => x"9387c4be",
        2273 => x"1304c4be",
        2274 => x"3304f440",
        2275 => x"13542440",
        2276 => x"9384c4be",
        2277 => x"13090000",
        2278 => x"63188902",
        2279 => x"8320c100",
        2280 => x"03248100",
        2281 => x"83244100",
        2282 => x"03290100",
        2283 => x"13010101",
        2284 => x"67800000",
        2285 => x"83a70400",
        2286 => x"13091900",
        2287 => x"93844400",
        2288 => x"e7800700",
        2289 => x"6ff01ffb",
        2290 => x"83a70400",
        2291 => x"13091900",
        2292 => x"93844400",
        2293 => x"e7800700",
        2294 => x"6ff01ffc",
        2295 => x"13860500",
        2296 => x"93050500",
        2297 => x"03a54187",
        2298 => x"6f10401e",
        2299 => x"638a050e",
        2300 => x"83a7c5ff",
        2301 => x"130101fe",
        2302 => x"232c8100",
        2303 => x"232e1100",
        2304 => x"1384c5ff",
        2305 => x"63d40700",
        2306 => x"3304f400",
        2307 => x"2326a100",
        2308 => x"ef008031",
        2309 => x"83a7c188",
        2310 => x"0325c100",
        2311 => x"639e0700",
        2312 => x"23220400",
        2313 => x"23a68188",
        2314 => x"03248101",
        2315 => x"8320c101",
        2316 => x"13010102",
        2317 => x"6f00802f",
        2318 => x"6374f402",
        2319 => x"03260400",
        2320 => x"b306c400",
        2321 => x"639ad700",
        2322 => x"83a60700",
        2323 => x"83a74700",
        2324 => x"b386c600",
        2325 => x"2320d400",
        2326 => x"2322f400",
        2327 => x"6ff09ffc",
        2328 => x"13870700",
        2329 => x"83a74700",
        2330 => x"63840700",
        2331 => x"e37af4fe",
        2332 => x"83260700",
        2333 => x"3306d700",
        2334 => x"63188602",
        2335 => x"03260400",
        2336 => x"b386c600",
        2337 => x"2320d700",
        2338 => x"3306d700",
        2339 => x"e39ec7f8",
        2340 => x"03a60700",
        2341 => x"83a74700",
        2342 => x"b306d600",
        2343 => x"2320d700",
        2344 => x"2322f700",
        2345 => x"6ff05ff8",
        2346 => x"6378c400",
        2347 => x"9307c000",
        2348 => x"2320f500",
        2349 => x"6ff05ff7",
        2350 => x"03260400",
        2351 => x"b306c400",
        2352 => x"639ad700",
        2353 => x"83a60700",
        2354 => x"83a74700",
        2355 => x"b386c600",
        2356 => x"2320d400",
        2357 => x"2322f400",
        2358 => x"23228700",
        2359 => x"6ff0dff4",
        2360 => x"67800000",
        2361 => x"130101ff",
        2362 => x"23202101",
        2363 => x"83a78188",
        2364 => x"23248100",
        2365 => x"23229100",
        2366 => x"23261100",
        2367 => x"93040500",
        2368 => x"13840500",
        2369 => x"63980700",
        2370 => x"93050000",
        2371 => x"ef10c010",
        2372 => x"23a4a188",
        2373 => x"93050400",
        2374 => x"13850400",
        2375 => x"ef10c00f",
        2376 => x"1309f0ff",
        2377 => x"63122503",
        2378 => x"1304f0ff",
        2379 => x"8320c100",
        2380 => x"13050400",
        2381 => x"03248100",
        2382 => x"83244100",
        2383 => x"03290100",
        2384 => x"13010101",
        2385 => x"67800000",
        2386 => x"13043500",
        2387 => x"1374c4ff",
        2388 => x"e30e85fc",
        2389 => x"b305a440",
        2390 => x"13850400",
        2391 => x"ef10c00b",
        2392 => x"e31625fd",
        2393 => x"6ff05ffc",
        2394 => x"130101fe",
        2395 => x"232a9100",
        2396 => x"93843500",
        2397 => x"93f4c4ff",
        2398 => x"23282101",
        2399 => x"232e1100",
        2400 => x"232c8100",
        2401 => x"23263101",
        2402 => x"23244101",
        2403 => x"93848400",
        2404 => x"9307c000",
        2405 => x"13090500",
        2406 => x"63f0f40a",
        2407 => x"9304c000",
        2408 => x"63eeb408",
        2409 => x"13050900",
        2410 => x"ef000018",
        2411 => x"83a7c188",
        2412 => x"13840700",
        2413 => x"631a040a",
        2414 => x"93850400",
        2415 => x"13050900",
        2416 => x"eff05ff2",
        2417 => x"9307f0ff",
        2418 => x"13040500",
        2419 => x"6316f514",
        2420 => x"03a4c188",
        2421 => x"93070400",
        2422 => x"639c0710",
        2423 => x"63040412",
        2424 => x"032a0400",
        2425 => x"93050000",
        2426 => x"13050900",
        2427 => x"330a4401",
        2428 => x"ef108002",
        2429 => x"6318aa10",
        2430 => x"83270400",
        2431 => x"13050900",
        2432 => x"b384f440",
        2433 => x"93850400",
        2434 => x"eff0dfed",
        2435 => x"9307f0ff",
        2436 => x"630af50e",
        2437 => x"83270400",
        2438 => x"b3879700",
        2439 => x"2320f400",
        2440 => x"83a7c188",
        2441 => x"638e070e",
        2442 => x"03a74700",
        2443 => x"6318870c",
        2444 => x"23a20700",
        2445 => x"6f004006",
        2446 => x"e3d404f6",
        2447 => x"9307c000",
        2448 => x"2320f900",
        2449 => x"13050000",
        2450 => x"8320c101",
        2451 => x"03248101",
        2452 => x"83244101",
        2453 => x"03290101",
        2454 => x"8329c100",
        2455 => x"032a8100",
        2456 => x"13010102",
        2457 => x"67800000",
        2458 => x"83260400",
        2459 => x"b3869640",
        2460 => x"63ca0606",
        2461 => x"1307b000",
        2462 => x"637ad704",
        2463 => x"23209400",
        2464 => x"33079400",
        2465 => x"63908704",
        2466 => x"23a6e188",
        2467 => x"83274400",
        2468 => x"2320d700",
        2469 => x"2322f700",
        2470 => x"13050900",
        2471 => x"ef000009",
        2472 => x"1305b400",
        2473 => x"93074400",
        2474 => x"137585ff",
        2475 => x"3307f540",
        2476 => x"e30cf5f8",
        2477 => x"3304e400",
        2478 => x"b387a740",
        2479 => x"2320f400",
        2480 => x"6ff09ff8",
        2481 => x"23a2e700",
        2482 => x"6ff05ffc",
        2483 => x"03274400",
        2484 => x"63968700",
        2485 => x"23a6e188",
        2486 => x"6ff01ffc",
        2487 => x"23a2e700",
        2488 => x"6ff09ffb",
        2489 => x"93070400",
        2490 => x"03244400",
        2491 => x"6ff09fec",
        2492 => x"13840700",
        2493 => x"83a74700",
        2494 => x"6ff01fee",
        2495 => x"93070700",
        2496 => x"6ff05ff2",
        2497 => x"9307c000",
        2498 => x"2320f900",
        2499 => x"13050900",
        2500 => x"ef00c001",
        2501 => x"6ff01ff3",
        2502 => x"23209500",
        2503 => x"6ff0dff7",
        2504 => x"23220000",
        2505 => x"73001000",
        2506 => x"67800000",
        2507 => x"67800000",
        2508 => x"130101fe",
        2509 => x"23282101",
        2510 => x"03a98500",
        2511 => x"232c8100",
        2512 => x"23263101",
        2513 => x"23225101",
        2514 => x"23206101",
        2515 => x"232e1100",
        2516 => x"232a9100",
        2517 => x"23244101",
        2518 => x"83aa0500",
        2519 => x"13840500",
        2520 => x"130b0600",
        2521 => x"93890600",
        2522 => x"63ec2609",
        2523 => x"8397c500",
        2524 => x"13f70748",
        2525 => x"63040708",
        2526 => x"03274401",
        2527 => x"93043000",
        2528 => x"83a50501",
        2529 => x"b384e402",
        2530 => x"13072000",
        2531 => x"b38aba40",
        2532 => x"130a0500",
        2533 => x"b3c4e402",
        2534 => x"13871600",
        2535 => x"33075701",
        2536 => x"63f4e400",
        2537 => x"93040700",
        2538 => x"93f70740",
        2539 => x"6386070a",
        2540 => x"93850400",
        2541 => x"13050a00",
        2542 => x"eff01fdb",
        2543 => x"13090500",
        2544 => x"630c050a",
        2545 => x"83250401",
        2546 => x"13860a00",
        2547 => x"efe01fbb",
        2548 => x"8357c400",
        2549 => x"93f7f7b7",
        2550 => x"93e70708",
        2551 => x"2316f400",
        2552 => x"23282401",
        2553 => x"232a9400",
        2554 => x"33095901",
        2555 => x"b3845441",
        2556 => x"23202401",
        2557 => x"23249400",
        2558 => x"13890900",
        2559 => x"63f42901",
        2560 => x"13890900",
        2561 => x"03250400",
        2562 => x"13060900",
        2563 => x"93050b00",
        2564 => x"efe01fb9",
        2565 => x"83278400",
        2566 => x"13050000",
        2567 => x"b3872741",
        2568 => x"2324f400",
        2569 => x"83270400",
        2570 => x"b3872701",
        2571 => x"2320f400",
        2572 => x"8320c101",
        2573 => x"03248101",
        2574 => x"83244101",
        2575 => x"03290101",
        2576 => x"8329c100",
        2577 => x"032a8100",
        2578 => x"832a4100",
        2579 => x"032b0100",
        2580 => x"13010102",
        2581 => x"67800000",
        2582 => x"13860400",
        2583 => x"13050a00",
        2584 => x"ef001060",
        2585 => x"13090500",
        2586 => x"e31c05f6",
        2587 => x"83250401",
        2588 => x"13050a00",
        2589 => x"eff09fb7",
        2590 => x"9307c000",
        2591 => x"2320fa00",
        2592 => x"8357c400",
        2593 => x"1305f0ff",
        2594 => x"93e70704",
        2595 => x"2316f400",
        2596 => x"6ff01ffa",
        2597 => x"83278600",
        2598 => x"130101fd",
        2599 => x"232e3101",
        2600 => x"23267101",
        2601 => x"23261102",
        2602 => x"23248102",
        2603 => x"23229102",
        2604 => x"23202103",
        2605 => x"232c4101",
        2606 => x"232a5101",
        2607 => x"23286101",
        2608 => x"23248101",
        2609 => x"23229101",
        2610 => x"2320a101",
        2611 => x"832b0600",
        2612 => x"93090600",
        2613 => x"63980712",
        2614 => x"13050000",
        2615 => x"8320c102",
        2616 => x"03248102",
        2617 => x"23a20900",
        2618 => x"83244102",
        2619 => x"03290102",
        2620 => x"8329c101",
        2621 => x"032a8101",
        2622 => x"832a4101",
        2623 => x"032b0101",
        2624 => x"832bc100",
        2625 => x"032c8100",
        2626 => x"832c4100",
        2627 => x"032d0100",
        2628 => x"13010103",
        2629 => x"67800000",
        2630 => x"03ab0b00",
        2631 => x"03ad4b00",
        2632 => x"938b8b00",
        2633 => x"03298400",
        2634 => x"832a0400",
        2635 => x"e3060dfe",
        2636 => x"63642d09",
        2637 => x"8317c400",
        2638 => x"13f70748",
        2639 => x"63020708",
        2640 => x"83244401",
        2641 => x"83250401",
        2642 => x"b3049c02",
        2643 => x"b38aba40",
        2644 => x"13871a00",
        2645 => x"3307a701",
        2646 => x"b3c49403",
        2647 => x"63f4e400",
        2648 => x"93040700",
        2649 => x"93f70740",
        2650 => x"638c070a",
        2651 => x"93850400",
        2652 => x"13050a00",
        2653 => x"eff05fbf",
        2654 => x"13090500",
        2655 => x"6302050c",
        2656 => x"83250401",
        2657 => x"13860a00",
        2658 => x"efe05f9f",
        2659 => x"8357c400",
        2660 => x"93f7f7b7",
        2661 => x"93e70708",
        2662 => x"2316f400",
        2663 => x"23282401",
        2664 => x"232a9400",
        2665 => x"33095901",
        2666 => x"b3845441",
        2667 => x"23202401",
        2668 => x"23249400",
        2669 => x"13090d00",
        2670 => x"63742d01",
        2671 => x"13090d00",
        2672 => x"03250400",
        2673 => x"93050b00",
        2674 => x"13060900",
        2675 => x"efe05f9d",
        2676 => x"83278400",
        2677 => x"330bab01",
        2678 => x"b3872741",
        2679 => x"2324f400",
        2680 => x"83270400",
        2681 => x"b3872701",
        2682 => x"2320f400",
        2683 => x"83a78900",
        2684 => x"b387a741",
        2685 => x"23a4f900",
        2686 => x"e38007ee",
        2687 => x"130d0000",
        2688 => x"6ff05ff2",
        2689 => x"130a0500",
        2690 => x"13840500",
        2691 => x"130b0000",
        2692 => x"130d0000",
        2693 => x"130c3000",
        2694 => x"930c2000",
        2695 => x"6ff09ff0",
        2696 => x"13860400",
        2697 => x"13050a00",
        2698 => x"ef009043",
        2699 => x"13090500",
        2700 => x"e31605f6",
        2701 => x"83250401",
        2702 => x"13050a00",
        2703 => x"eff01f9b",
        2704 => x"9307c000",
        2705 => x"2320fa00",
        2706 => x"8357c400",
        2707 => x"1305f0ff",
        2708 => x"93e70704",
        2709 => x"2316f400",
        2710 => x"23a40900",
        2711 => x"6ff01fe8",
        2712 => x"83d7c500",
        2713 => x"130101f5",
        2714 => x"2324810a",
        2715 => x"2322910a",
        2716 => x"2320210b",
        2717 => x"232c4109",
        2718 => x"2326110a",
        2719 => x"232e3109",
        2720 => x"232a5109",
        2721 => x"23286109",
        2722 => x"23267109",
        2723 => x"23248109",
        2724 => x"23229109",
        2725 => x"2320a109",
        2726 => x"232eb107",
        2727 => x"93f70708",
        2728 => x"130a0500",
        2729 => x"13890500",
        2730 => x"93040600",
        2731 => x"13840600",
        2732 => x"63880706",
        2733 => x"83a70501",
        2734 => x"63940706",
        2735 => x"93050004",
        2736 => x"eff09faa",
        2737 => x"2320a900",
        2738 => x"2328a900",
        2739 => x"63160504",
        2740 => x"9307c000",
        2741 => x"2320fa00",
        2742 => x"1305f0ff",
        2743 => x"8320c10a",
        2744 => x"0324810a",
        2745 => x"8324410a",
        2746 => x"0329010a",
        2747 => x"8329c109",
        2748 => x"032a8109",
        2749 => x"832a4109",
        2750 => x"032b0109",
        2751 => x"832bc108",
        2752 => x"032c8108",
        2753 => x"832c4108",
        2754 => x"032d0108",
        2755 => x"832dc107",
        2756 => x"1301010b",
        2757 => x"67800000",
        2758 => x"93070004",
        2759 => x"232af900",
        2760 => x"93070002",
        2761 => x"a304f102",
        2762 => x"93070003",
        2763 => x"23220102",
        2764 => x"2305f102",
        2765 => x"23268100",
        2766 => x"930c5002",
        2767 => x"374b0000",
        2768 => x"b74b0000",
        2769 => x"374d0000",
        2770 => x"372c0000",
        2771 => x"930a0000",
        2772 => x"13840400",
        2773 => x"83470400",
        2774 => x"63840700",
        2775 => x"639c970d",
        2776 => x"b30d9440",
        2777 => x"63069402",
        2778 => x"93860d00",
        2779 => x"13860400",
        2780 => x"93050900",
        2781 => x"13050a00",
        2782 => x"eff09fbb",
        2783 => x"9307f0ff",
        2784 => x"6304f524",
        2785 => x"83274102",
        2786 => x"b387b701",
        2787 => x"2322f102",
        2788 => x"83470400",
        2789 => x"638a0722",
        2790 => x"9307f0ff",
        2791 => x"93041400",
        2792 => x"23280100",
        2793 => x"232e0100",
        2794 => x"232af100",
        2795 => x"232c0100",
        2796 => x"a3090104",
        2797 => x"23240106",
        2798 => x"930d1000",
        2799 => x"83c50400",
        2800 => x"13065000",
        2801 => x"13058bb5",
        2802 => x"ef00101e",
        2803 => x"83270101",
        2804 => x"13841400",
        2805 => x"63140506",
        2806 => x"13f70701",
        2807 => x"63060700",
        2808 => x"13070002",
        2809 => x"a309e104",
        2810 => x"13f78700",
        2811 => x"63060700",
        2812 => x"1307b002",
        2813 => x"a309e104",
        2814 => x"83c60400",
        2815 => x"1307a002",
        2816 => x"638ce604",
        2817 => x"8327c101",
        2818 => x"13840400",
        2819 => x"93060000",
        2820 => x"13069000",
        2821 => x"1305a000",
        2822 => x"03470400",
        2823 => x"93051400",
        2824 => x"130707fd",
        2825 => x"637ee608",
        2826 => x"63840604",
        2827 => x"232ef100",
        2828 => x"6f000004",
        2829 => x"13041400",
        2830 => x"6ff0dff1",
        2831 => x"13078bb5",
        2832 => x"3305e540",
        2833 => x"3395ad00",
        2834 => x"b3e7a700",
        2835 => x"2328f100",
        2836 => x"93040400",
        2837 => x"6ff09ff6",
        2838 => x"0327c100",
        2839 => x"93064700",
        2840 => x"03270700",
        2841 => x"2326d100",
        2842 => x"63420704",
        2843 => x"232ee100",
        2844 => x"03470400",
        2845 => x"9307e002",
        2846 => x"6314f708",
        2847 => x"03471400",
        2848 => x"9307a002",
        2849 => x"6318f704",
        2850 => x"8327c100",
        2851 => x"13042400",
        2852 => x"13874700",
        2853 => x"83a70700",
        2854 => x"2326e100",
        2855 => x"63d40700",
        2856 => x"9307f0ff",
        2857 => x"232af100",
        2858 => x"6f008005",
        2859 => x"3307e040",
        2860 => x"93e72700",
        2861 => x"232ee100",
        2862 => x"2328f100",
        2863 => x"6ff05ffb",
        2864 => x"b387a702",
        2865 => x"13840500",
        2866 => x"93061000",
        2867 => x"b387e700",
        2868 => x"6ff09ff4",
        2869 => x"13041400",
        2870 => x"232a0100",
        2871 => x"93060000",
        2872 => x"93070000",
        2873 => x"13069000",
        2874 => x"1305a000",
        2875 => x"03470400",
        2876 => x"93051400",
        2877 => x"130707fd",
        2878 => x"6372e608",
        2879 => x"e39406fa",
        2880 => x"83450400",
        2881 => x"13063000",
        2882 => x"13850bb6",
        2883 => x"ef00d009",
        2884 => x"63020502",
        2885 => x"93870bb6",
        2886 => x"3305f540",
        2887 => x"83270101",
        2888 => x"13070004",
        2889 => x"3317a700",
        2890 => x"b3e7e700",
        2891 => x"13041400",
        2892 => x"2328f100",
        2893 => x"83450400",
        2894 => x"13066000",
        2895 => x"13054db6",
        2896 => x"93041400",
        2897 => x"2304b102",
        2898 => x"ef001006",
        2899 => x"63080508",
        2900 => x"63980a04",
        2901 => x"03270101",
        2902 => x"8327c100",
        2903 => x"13770710",
        2904 => x"63080702",
        2905 => x"93874700",
        2906 => x"2326f100",
        2907 => x"83274102",
        2908 => x"b3873701",
        2909 => x"2322f102",
        2910 => x"6ff09fdd",
        2911 => x"b387a702",
        2912 => x"13840500",
        2913 => x"93061000",
        2914 => x"b387e700",
        2915 => x"6ff01ff6",
        2916 => x"93877700",
        2917 => x"93f787ff",
        2918 => x"93878700",
        2919 => x"6ff0dffc",
        2920 => x"1307c100",
        2921 => x"93060c73",
        2922 => x"13060900",
        2923 => x"93050101",
        2924 => x"13050a00",
        2925 => x"97000000",
        2926 => x"e7000000",
        2927 => x"9307f0ff",
        2928 => x"93090500",
        2929 => x"e314f5fa",
        2930 => x"8357c900",
        2931 => x"93f70704",
        2932 => x"e39407d0",
        2933 => x"03254102",
        2934 => x"6ff05fd0",
        2935 => x"1307c100",
        2936 => x"93060c73",
        2937 => x"13060900",
        2938 => x"93050101",
        2939 => x"13050a00",
        2940 => x"ef00801b",
        2941 => x"6ff09ffc",
        2942 => x"130101fd",
        2943 => x"232a5101",
        2944 => x"83a70501",
        2945 => x"930a0700",
        2946 => x"03a78500",
        2947 => x"23248102",
        2948 => x"23202103",
        2949 => x"232e3101",
        2950 => x"232c4101",
        2951 => x"23261102",
        2952 => x"23229102",
        2953 => x"23286101",
        2954 => x"23267101",
        2955 => x"93090500",
        2956 => x"13840500",
        2957 => x"13090600",
        2958 => x"138a0600",
        2959 => x"63d4e700",
        2960 => x"93070700",
        2961 => x"2320f900",
        2962 => x"03473404",
        2963 => x"63060700",
        2964 => x"93871700",
        2965 => x"2320f900",
        2966 => x"83270400",
        2967 => x"93f70702",
        2968 => x"63880700",
        2969 => x"83270900",
        2970 => x"93872700",
        2971 => x"2320f900",
        2972 => x"83240400",
        2973 => x"93f46400",
        2974 => x"639e0400",
        2975 => x"130b9401",
        2976 => x"930bf0ff",
        2977 => x"8327c400",
        2978 => x"03270900",
        2979 => x"b387e740",
        2980 => x"63c2f408",
        2981 => x"83473404",
        2982 => x"b336f000",
        2983 => x"83270400",
        2984 => x"93f70702",
        2985 => x"6390070c",
        2986 => x"13063404",
        2987 => x"93050a00",
        2988 => x"13850900",
        2989 => x"e7800a00",
        2990 => x"9307f0ff",
        2991 => x"6308f506",
        2992 => x"83270400",
        2993 => x"13074000",
        2994 => x"93040000",
        2995 => x"93f76700",
        2996 => x"639ce700",
        2997 => x"8324c400",
        2998 => x"83270900",
        2999 => x"b384f440",
        3000 => x"63d40400",
        3001 => x"93040000",
        3002 => x"83278400",
        3003 => x"03270401",
        3004 => x"6356f700",
        3005 => x"b387e740",
        3006 => x"b384f400",
        3007 => x"13090000",
        3008 => x"1304a401",
        3009 => x"130bf0ff",
        3010 => x"63902409",
        3011 => x"13050000",
        3012 => x"6f000002",
        3013 => x"93061000",
        3014 => x"13060b00",
        3015 => x"93050a00",
        3016 => x"13850900",
        3017 => x"e7800a00",
        3018 => x"631a7503",
        3019 => x"1305f0ff",
        3020 => x"8320c102",
        3021 => x"03248102",
        3022 => x"83244102",
        3023 => x"03290102",
        3024 => x"8329c101",
        3025 => x"032a8101",
        3026 => x"832a4101",
        3027 => x"032b0101",
        3028 => x"832bc100",
        3029 => x"13010103",
        3030 => x"67800000",
        3031 => x"93841400",
        3032 => x"6ff05ff2",
        3033 => x"3307d400",
        3034 => x"13060003",
        3035 => x"a301c704",
        3036 => x"03475404",
        3037 => x"93871600",
        3038 => x"b307f400",
        3039 => x"93862600",
        3040 => x"a381e704",
        3041 => x"6ff05ff2",
        3042 => x"93061000",
        3043 => x"13060400",
        3044 => x"93050a00",
        3045 => x"13850900",
        3046 => x"e7800a00",
        3047 => x"e30865f9",
        3048 => x"13091900",
        3049 => x"6ff05ff6",
        3050 => x"130101fd",
        3051 => x"23248102",
        3052 => x"23202103",
        3053 => x"232e3101",
        3054 => x"232c4101",
        3055 => x"23261102",
        3056 => x"23229102",
        3057 => x"232a5101",
        3058 => x"23286101",
        3059 => x"138a0600",
        3060 => x"83c68501",
        3061 => x"93078007",
        3062 => x"13090500",
        3063 => x"13840500",
        3064 => x"93090600",
        3065 => x"63eed700",
        3066 => x"93072006",
        3067 => x"13863504",
        3068 => x"63eed700",
        3069 => x"63840628",
        3070 => x"93078005",
        3071 => x"6380f622",
        3072 => x"93042404",
        3073 => x"2301d404",
        3074 => x"6f004004",
        3075 => x"9387d6f9",
        3076 => x"93f7f70f",
        3077 => x"93055001",
        3078 => x"e3e4f5fe",
        3079 => x"b7450000",
        3080 => x"93972700",
        3081 => x"938545b9",
        3082 => x"b387b700",
        3083 => x"83a70700",
        3084 => x"67800700",
        3085 => x"83270700",
        3086 => x"93042404",
        3087 => x"93864700",
        3088 => x"83a70700",
        3089 => x"2320d700",
        3090 => x"2301f404",
        3091 => x"93071000",
        3092 => x"6f008026",
        3093 => x"83270400",
        3094 => x"03250700",
        3095 => x"93f60708",
        3096 => x"93054500",
        3097 => x"63860602",
        3098 => x"83270500",
        3099 => x"2320b700",
        3100 => x"37480000",
        3101 => x"63d80700",
        3102 => x"1307d002",
        3103 => x"b307f040",
        3104 => x"a301e404",
        3105 => x"1308c8b6",
        3106 => x"1307a000",
        3107 => x"6f004006",
        3108 => x"93f60704",
        3109 => x"83270500",
        3110 => x"2320b700",
        3111 => x"e38a06fc",
        3112 => x"93970701",
        3113 => x"93d70741",
        3114 => x"6ff09ffc",
        3115 => x"03250400",
        3116 => x"83250700",
        3117 => x"13780508",
        3118 => x"83a70500",
        3119 => x"93854500",
        3120 => x"631a0800",
        3121 => x"13750504",
        3122 => x"63060500",
        3123 => x"93970701",
        3124 => x"93d70701",
        3125 => x"2320b700",
        3126 => x"37480000",
        3127 => x"1307f006",
        3128 => x"1308c8b6",
        3129 => x"639ae614",
        3130 => x"13078000",
        3131 => x"a3010404",
        3132 => x"83264400",
        3133 => x"2324d400",
        3134 => x"63ce0600",
        3135 => x"83250400",
        3136 => x"b3e6d700",
        3137 => x"93040600",
        3138 => x"93f5b5ff",
        3139 => x"2320b400",
        3140 => x"63840602",
        3141 => x"93040600",
        3142 => x"b3f6e702",
        3143 => x"9384f4ff",
        3144 => x"b306d800",
        3145 => x"83c60600",
        3146 => x"2380d400",
        3147 => x"93860700",
        3148 => x"b3d7e702",
        3149 => x"e3f2e6fe",
        3150 => x"93078000",
        3151 => x"6314f702",
        3152 => x"83270400",
        3153 => x"93f71700",
        3154 => x"638e0700",
        3155 => x"03274400",
        3156 => x"83270401",
        3157 => x"63c8e700",
        3158 => x"93070003",
        3159 => x"a38ff4fe",
        3160 => x"9384f4ff",
        3161 => x"33069640",
        3162 => x"2328c400",
        3163 => x"13070a00",
        3164 => x"93860900",
        3165 => x"1306c100",
        3166 => x"93050400",
        3167 => x"13050900",
        3168 => x"eff09fc7",
        3169 => x"930af0ff",
        3170 => x"631e5513",
        3171 => x"1305f0ff",
        3172 => x"8320c102",
        3173 => x"03248102",
        3174 => x"83244102",
        3175 => x"03290102",
        3176 => x"8329c101",
        3177 => x"032a8101",
        3178 => x"832a4101",
        3179 => x"032b0101",
        3180 => x"13010103",
        3181 => x"67800000",
        3182 => x"83270400",
        3183 => x"93e70702",
        3184 => x"2320f400",
        3185 => x"37480000",
        3186 => x"93068007",
        3187 => x"130808b8",
        3188 => x"a302d404",
        3189 => x"83260400",
        3190 => x"83250700",
        3191 => x"13f50608",
        3192 => x"83a70500",
        3193 => x"93854500",
        3194 => x"631a0500",
        3195 => x"13f50604",
        3196 => x"63060500",
        3197 => x"93970701",
        3198 => x"93d70701",
        3199 => x"2320b700",
        3200 => x"13f71600",
        3201 => x"63060700",
        3202 => x"93e60602",
        3203 => x"2320d400",
        3204 => x"638c0700",
        3205 => x"13070001",
        3206 => x"6ff05fed",
        3207 => x"37480000",
        3208 => x"1308c8b6",
        3209 => x"6ff0dffa",
        3210 => x"03270400",
        3211 => x"1377f7fd",
        3212 => x"2320e400",
        3213 => x"6ff01ffe",
        3214 => x"1307a000",
        3215 => x"6ff01feb",
        3216 => x"83260400",
        3217 => x"83270700",
        3218 => x"83254401",
        3219 => x"13f80608",
        3220 => x"13854700",
        3221 => x"630a0800",
        3222 => x"2320a700",
        3223 => x"83a70700",
        3224 => x"23a0b700",
        3225 => x"6f008001",
        3226 => x"2320a700",
        3227 => x"93f60604",
        3228 => x"83a70700",
        3229 => x"e38606fe",
        3230 => x"2390b700",
        3231 => x"23280400",
        3232 => x"93040600",
        3233 => x"6ff09fee",
        3234 => x"83270700",
        3235 => x"03264400",
        3236 => x"93050000",
        3237 => x"93864700",
        3238 => x"2320d700",
        3239 => x"83a40700",
        3240 => x"13850400",
        3241 => x"ef004030",
        3242 => x"63060500",
        3243 => x"33059540",
        3244 => x"2322a400",
        3245 => x"83274400",
        3246 => x"2328f400",
        3247 => x"a3010404",
        3248 => x"6ff0dfea",
        3249 => x"83260401",
        3250 => x"13860400",
        3251 => x"93850900",
        3252 => x"13050900",
        3253 => x"e7000a00",
        3254 => x"e30a55eb",
        3255 => x"83270400",
        3256 => x"93f72700",
        3257 => x"63940704",
        3258 => x"8327c100",
        3259 => x"0325c400",
        3260 => x"e350f5ea",
        3261 => x"13850700",
        3262 => x"6ff09fe9",
        3263 => x"93061000",
        3264 => x"13860a00",
        3265 => x"93850900",
        3266 => x"13050900",
        3267 => x"e7000a00",
        3268 => x"e30e65e7",
        3269 => x"93841400",
        3270 => x"8327c400",
        3271 => x"0327c100",
        3272 => x"b387e740",
        3273 => x"e3ccf4fc",
        3274 => x"6ff01ffc",
        3275 => x"93040000",
        3276 => x"930a9401",
        3277 => x"130bf0ff",
        3278 => x"6ff01ffe",
        3279 => x"8397c500",
        3280 => x"130101fe",
        3281 => x"232c8100",
        3282 => x"232a9100",
        3283 => x"232e1100",
        3284 => x"23282101",
        3285 => x"23263101",
        3286 => x"13f78700",
        3287 => x"93040500",
        3288 => x"13840500",
        3289 => x"631a0712",
        3290 => x"03a74500",
        3291 => x"6346e000",
        3292 => x"03a70504",
        3293 => x"6356e010",
        3294 => x"0327c402",
        3295 => x"63020710",
        3296 => x"03a90400",
        3297 => x"93963701",
        3298 => x"23a00400",
        3299 => x"83250402",
        3300 => x"63dc060a",
        3301 => x"03264405",
        3302 => x"8357c400",
        3303 => x"93f74700",
        3304 => x"638e0700",
        3305 => x"83274400",
        3306 => x"3306f640",
        3307 => x"83274403",
        3308 => x"63860700",
        3309 => x"83270404",
        3310 => x"3306f640",
        3311 => x"8327c402",
        3312 => x"83250402",
        3313 => x"93060000",
        3314 => x"13850400",
        3315 => x"e7800700",
        3316 => x"1307f0ff",
        3317 => x"8357c400",
        3318 => x"6312e502",
        3319 => x"83a60400",
        3320 => x"1307d001",
        3321 => x"6362d70a",
        3322 => x"37074020",
        3323 => x"13071700",
        3324 => x"3357d700",
        3325 => x"13771700",
        3326 => x"63080708",
        3327 => x"03270401",
        3328 => x"23220400",
        3329 => x"2320e400",
        3330 => x"13973701",
        3331 => x"635c0700",
        3332 => x"9307f0ff",
        3333 => x"6316f500",
        3334 => x"83a70400",
        3335 => x"63940700",
        3336 => x"232aa404",
        3337 => x"83254403",
        3338 => x"23a02401",
        3339 => x"638a0504",
        3340 => x"93074404",
        3341 => x"6386f500",
        3342 => x"13850400",
        3343 => x"efe01ffb",
        3344 => x"232a0402",
        3345 => x"6f00c003",
        3346 => x"13060000",
        3347 => x"93061000",
        3348 => x"13850400",
        3349 => x"e7000700",
        3350 => x"9307f0ff",
        3351 => x"13060500",
        3352 => x"e31cf5f2",
        3353 => x"83a70400",
        3354 => x"e38807f2",
        3355 => x"1307d001",
        3356 => x"6386e700",
        3357 => x"13076001",
        3358 => x"6394e706",
        3359 => x"23a02401",
        3360 => x"13050000",
        3361 => x"6f00c006",
        3362 => x"93e70704",
        3363 => x"93970701",
        3364 => x"93d70741",
        3365 => x"6f004005",
        3366 => x"83a90501",
        3367 => x"e38209fe",
        3368 => x"03a90500",
        3369 => x"93f73700",
        3370 => x"23a03501",
        3371 => x"33093941",
        3372 => x"13070000",
        3373 => x"63940700",
        3374 => x"03a74501",
        3375 => x"2324e400",
        3376 => x"e35020fd",
        3377 => x"83278402",
        3378 => x"83250402",
        3379 => x"93060900",
        3380 => x"13860900",
        3381 => x"13850400",
        3382 => x"e7800700",
        3383 => x"6348a002",
        3384 => x"8317c400",
        3385 => x"93e70704",
        3386 => x"2316f400",
        3387 => x"1305f0ff",
        3388 => x"8320c101",
        3389 => x"03248101",
        3390 => x"83244101",
        3391 => x"03290101",
        3392 => x"8329c100",
        3393 => x"13010102",
        3394 => x"67800000",
        3395 => x"b389a900",
        3396 => x"3309a940",
        3397 => x"6ff0dffa",
        3398 => x"83a70501",
        3399 => x"638e0704",
        3400 => x"130101fe",
        3401 => x"232c8100",
        3402 => x"232e1100",
        3403 => x"13040500",
        3404 => x"630c0500",
        3405 => x"83270502",
        3406 => x"63980700",
        3407 => x"2326b100",
        3408 => x"efe05f85",
        3409 => x"8325c100",
        3410 => x"8397c500",
        3411 => x"638c0700",
        3412 => x"13050400",
        3413 => x"03248101",
        3414 => x"8320c101",
        3415 => x"13010102",
        3416 => x"6ff0dfdd",
        3417 => x"8320c101",
        3418 => x"03248101",
        3419 => x"13050000",
        3420 => x"13010102",
        3421 => x"67800000",
        3422 => x"13050000",
        3423 => x"67800000",
        3424 => x"93050500",
        3425 => x"631e0500",
        3426 => x"b7350000",
        3427 => x"37050020",
        3428 => x"13868181",
        3429 => x"93858551",
        3430 => x"13054502",
        3431 => x"6fe0df84",
        3432 => x"03a54187",
        3433 => x"6ff05ff7",
        3434 => x"93f5f50f",
        3435 => x"3306c500",
        3436 => x"6316c500",
        3437 => x"13050000",
        3438 => x"67800000",
        3439 => x"83470500",
        3440 => x"e38cb7fe",
        3441 => x"13051500",
        3442 => x"6ff09ffe",
        3443 => x"130101ff",
        3444 => x"23248100",
        3445 => x"23229100",
        3446 => x"13040500",
        3447 => x"13850500",
        3448 => x"93050600",
        3449 => x"23261100",
        3450 => x"23a20188",
        3451 => x"efd05fdf",
        3452 => x"9307f0ff",
        3453 => x"6318f500",
        3454 => x"83a74188",
        3455 => x"63840700",
        3456 => x"2320f400",
        3457 => x"8320c100",
        3458 => x"03248100",
        3459 => x"83244100",
        3460 => x"13010101",
        3461 => x"67800000",
        3462 => x"130101ff",
        3463 => x"23248100",
        3464 => x"23229100",
        3465 => x"13040500",
        3466 => x"13850500",
        3467 => x"23261100",
        3468 => x"23a20188",
        3469 => x"efe08f82",
        3470 => x"9307f0ff",
        3471 => x"6318f500",
        3472 => x"83a74188",
        3473 => x"63840700",
        3474 => x"2320f400",
        3475 => x"8320c100",
        3476 => x"03248100",
        3477 => x"83244100",
        3478 => x"13010101",
        3479 => x"67800000",
        3480 => x"130101fe",
        3481 => x"232c8100",
        3482 => x"232e1100",
        3483 => x"232a9100",
        3484 => x"23282101",
        3485 => x"23263101",
        3486 => x"23244101",
        3487 => x"13040600",
        3488 => x"63940502",
        3489 => x"03248101",
        3490 => x"8320c101",
        3491 => x"83244101",
        3492 => x"03290101",
        3493 => x"8329c100",
        3494 => x"032a8100",
        3495 => x"93050600",
        3496 => x"13010102",
        3497 => x"6fe05fec",
        3498 => x"63180602",
        3499 => x"efe01fd4",
        3500 => x"93040000",
        3501 => x"8320c101",
        3502 => x"03248101",
        3503 => x"03290101",
        3504 => x"8329c100",
        3505 => x"032a8100",
        3506 => x"13850400",
        3507 => x"83244101",
        3508 => x"13010102",
        3509 => x"67800000",
        3510 => x"130a0500",
        3511 => x"93840500",
        3512 => x"ef008005",
        3513 => x"13090500",
        3514 => x"63668500",
        3515 => x"93571500",
        3516 => x"e3e287fc",
        3517 => x"93050400",
        3518 => x"13050a00",
        3519 => x"efe0dfe6",
        3520 => x"93090500",
        3521 => x"63160500",
        3522 => x"93840900",
        3523 => x"6ff09ffa",
        3524 => x"13060400",
        3525 => x"63748900",
        3526 => x"13060900",
        3527 => x"93850400",
        3528 => x"13850900",
        3529 => x"efd09fc5",
        3530 => x"93850400",
        3531 => x"13050a00",
        3532 => x"efe0dfcb",
        3533 => x"6ff05ffd",
        3534 => x"83a7c5ff",
        3535 => x"1385c7ff",
        3536 => x"63d80700",
        3537 => x"b385a500",
        3538 => x"83a70500",
        3539 => x"3305f500",
        3540 => x"67800000",
        3541 => x"10000000",
        3542 => x"00000000",
        3543 => x"037a5200",
        3544 => x"017c0101",
        3545 => x"1b0d0200",
        3546 => x"10000000",
        3547 => x"18000000",
        3548 => x"64cfffff",
        3549 => x"78040000",
        3550 => x"00000000",
        3551 => x"10000000",
        3552 => x"00000000",
        3553 => x"037a5200",
        3554 => x"017c0101",
        3555 => x"1b0d0200",
        3556 => x"10000000",
        3557 => x"18000000",
        3558 => x"b4d3ffff",
        3559 => x"30040000",
        3560 => x"00000000",
        3561 => x"10000000",
        3562 => x"00000000",
        3563 => x"037a5200",
        3564 => x"017c0101",
        3565 => x"1b0d0200",
        3566 => x"10000000",
        3567 => x"18000000",
        3568 => x"bcd7ffff",
        3569 => x"e4030000",
        3570 => x"00000000",
        3571 => x"30313233",
        3572 => x"34353637",
        3573 => x"38396162",
        3574 => x"63646566",
        3575 => x"00000000",
        3576 => x"88040000",
        3577 => x"c0030000",
        3578 => x"c0030000",
        3579 => x"c0030000",
        3580 => x"c0030000",
        3581 => x"c0030000",
        3582 => x"c0030000",
        3583 => x"c0030000",
        3584 => x"c0030000",
        3585 => x"c0030000",
        3586 => x"c0030000",
        3587 => x"94040000",
        3588 => x"c0030000",
        3589 => x"a0040000",
        3590 => x"ac040000",
        3591 => x"c0030000",
        3592 => x"b8040000",
        3593 => x"c4040000",
        3594 => x"c0030000",
        3595 => x"d0040000",
        3596 => x"7c040000",
        3597 => x"c0030000",
        3598 => x"c0030000",
        3599 => x"c0030000",
        3600 => x"dc040000",
        3601 => x"c0030000",
        3602 => x"c0030000",
        3603 => x"c0030000",
        3604 => x"c0030000",
        3605 => x"c0030000",
        3606 => x"c0030000",
        3607 => x"c0030000",
        3608 => x"ec040000",
        3609 => x"80050000",
        3610 => x"98050000",
        3611 => x"c8050000",
        3612 => x"48050000",
        3613 => x"48050000",
        3614 => x"48050000",
        3615 => x"48050000",
        3616 => x"48050000",
        3617 => x"48050000",
        3618 => x"b0050000",
        3619 => x"48050000",
        3620 => x"48050000",
        3621 => x"48050000",
        3622 => x"48050000",
        3623 => x"60050000",
        3624 => x"60050000",
        3625 => x"80050000",
        3626 => x"48050000",
        3627 => x"48050000",
        3628 => x"48050000",
        3629 => x"48050000",
        3630 => x"74050000",
        3631 => x"e0050000",
        3632 => x"08060000",
        3633 => x"48050000",
        3634 => x"48050000",
        3635 => x"48050000",
        3636 => x"48050000",
        3637 => x"48050000",
        3638 => x"48050000",
        3639 => x"48050000",
        3640 => x"48050000",
        3641 => x"48050000",
        3642 => x"48050000",
        3643 => x"48050000",
        3644 => x"48050000",
        3645 => x"48050000",
        3646 => x"48050000",
        3647 => x"60050000",
        3648 => x"60050000",
        3649 => x"48050000",
        3650 => x"48050000",
        3651 => x"48050000",
        3652 => x"48050000",
        3653 => x"48050000",
        3654 => x"48050000",
        3655 => x"48050000",
        3656 => x"48050000",
        3657 => x"48050000",
        3658 => x"48050000",
        3659 => x"48050000",
        3660 => x"48050000",
        3661 => x"74050000",
        3662 => x"00010202",
        3663 => x"03030303",
        3664 => x"04040404",
        3665 => x"04040404",
        3666 => x"05050505",
        3667 => x"05050505",
        3668 => x"05050505",
        3669 => x"05050505",
        3670 => x"06060606",
        3671 => x"06060606",
        3672 => x"06060606",
        3673 => x"06060606",
        3674 => x"06060606",
        3675 => x"06060606",
        3676 => x"06060606",
        3677 => x"06060606",
        3678 => x"07070707",
        3679 => x"07070707",
        3680 => x"07070707",
        3681 => x"07070707",
        3682 => x"07070707",
        3683 => x"07070707",
        3684 => x"07070707",
        3685 => x"07070707",
        3686 => x"07070707",
        3687 => x"07070707",
        3688 => x"07070707",
        3689 => x"07070707",
        3690 => x"07070707",
        3691 => x"07070707",
        3692 => x"07070707",
        3693 => x"07070707",
        3694 => x"08080808",
        3695 => x"08080808",
        3696 => x"08080808",
        3697 => x"08080808",
        3698 => x"08080808",
        3699 => x"08080808",
        3700 => x"08080808",
        3701 => x"08080808",
        3702 => x"08080808",
        3703 => x"08080808",
        3704 => x"08080808",
        3705 => x"08080808",
        3706 => x"08080808",
        3707 => x"08080808",
        3708 => x"08080808",
        3709 => x"08080808",
        3710 => x"08080808",
        3711 => x"08080808",
        3712 => x"08080808",
        3713 => x"08080808",
        3714 => x"08080808",
        3715 => x"08080808",
        3716 => x"08080808",
        3717 => x"08080808",
        3718 => x"08080808",
        3719 => x"08080808",
        3720 => x"08080808",
        3721 => x"08080808",
        3722 => x"08080808",
        3723 => x"08080808",
        3724 => x"08080808",
        3725 => x"08080808",
        3726 => x"0d0a4542",
        3727 => x"5245414b",
        3728 => x"21206d65",
        3729 => x"7063203d",
        3730 => x"20000000",
        3731 => x"20696e73",
        3732 => x"6e203d20",
        3733 => x"00000000",
        3734 => x"0d0a0000",
        3735 => x"0d0a0a44",
        3736 => x"6973706c",
        3737 => x"6179696e",
        3738 => x"67207468",
        3739 => x"65207469",
        3740 => x"6d652070",
        3741 => x"61737365",
        3742 => x"64207369",
        3743 => x"6e636520",
        3744 => x"72657365",
        3745 => x"740d0a0a",
        3746 => x"00000000",
        3747 => x"2530356c",
        3748 => x"643a2530",
        3749 => x"366c6420",
        3750 => x"20202530",
        3751 => x"326c643a",
        3752 => x"2530326c",
        3753 => x"643a2530",
        3754 => x"326c640d",
        3755 => x"00000000",
        3756 => x"696e7465",
        3757 => x"72727570",
        3758 => x"745f6469",
        3759 => x"72656374",
        3760 => x"00000000",
        3761 => x"54485541",
        3762 => x"53205249",
        3763 => x"53432d56",
        3764 => x"20525633",
        3765 => x"32494d20",
        3766 => x"62617265",
        3767 => x"206d6574",
        3768 => x"616c2070",
        3769 => x"726f6365",
        3770 => x"73736f72",
        3771 => x"00000000",
        3772 => x"54686520",
        3773 => x"48616775",
        3774 => x"6520556e",
        3775 => x"69766572",
        3776 => x"73697479",
        3777 => x"206f6620",
        3778 => x"4170706c",
        3779 => x"69656420",
        3780 => x"53636965",
        3781 => x"6e636573",
        3782 => x"00000000",
        3783 => x"44657061",
        3784 => x"72746d65",
        3785 => x"6e74206f",
        3786 => x"6620456c",
        3787 => x"65637472",
        3788 => x"6963616c",
        3789 => x"20456e67",
        3790 => x"696e6565",
        3791 => x"72696e67",
        3792 => x"00000000",
        3793 => x"4a2e452e",
        3794 => x"4a2e206f",
        3795 => x"70206465",
        3796 => x"6e204272",
        3797 => x"6f757700",
        3798 => x"232d302b",
        3799 => x"20000000",
        3800 => x"686c4c00",
        3801 => x"65666745",
        3802 => x"46470000",
        3803 => x"30313233",
        3804 => x"34353637",
        3805 => x"38394142",
        3806 => x"43444546",
        3807 => x"00000000",
        3808 => x"30313233",
        3809 => x"34353637",
        3810 => x"38396162",
        3811 => x"63646566",
        3812 => x"00000000",
        3813 => x"34300000",
        3814 => x"54300000",
        3815 => x"00300000",
        3816 => x"00300000",
        3817 => x"00300000",
        3818 => x"00300000",
        3819 => x"54300000",
        3820 => x"00300000",
        3821 => x"00300000",
        3822 => x"00300000",
        3823 => x"00300000",
        3824 => x"40320000",
        3825 => x"ac300000",
        3826 => x"b8310000",
        3827 => x"00300000",
        3828 => x"00300000",
        3829 => x"88320000",
        3830 => x"00300000",
        3831 => x"ac300000",
        3832 => x"00300000",
        3833 => x"00300000",
        3834 => x"c4310000",
        3835 => x"b03a0000",
        3836 => x"c43a0000",
        3837 => x"f03a0000",
        3838 => x"1c3b0000",
        3839 => x"443b0000",
        3840 => x"00000000",
        3841 => x"00000000",
        3842 => x"03000000",
        3843 => x"90000020",
        3844 => x"00000000",
        3845 => x"90000020",
        3846 => x"f8000020",
        3847 => x"60010020",
        3848 => x"00000000",
        3849 => x"00000000",
        3850 => x"00000000",
        3851 => x"00000000",
        3852 => x"00000000",
        3853 => x"00000000",
        3854 => x"00000000",
        3855 => x"00000000",
        3856 => x"00000000",
        3857 => x"00000000",
        3858 => x"00000000",
        3859 => x"00000000",
        3860 => x"00000000",
        3861 => x"00000000",
        3862 => x"00000000",
        3863 => x"78000020",
        3864 => x"24000020"
            );
end package rom_image;
