-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Thu Oct 19 19:01:28 2023


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382022b",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"13868187",
           8 => x"9387819c",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13858187",
          13 => x"ef10c02f",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93878187",
          17 => x"637cf600",
          18 => x"b7450000",
          19 => x"3386c740",
          20 => x"938585b6",
          21 => x"13050500",
          22 => x"ef10402f",
          23 => x"ef20c027",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10006d",
          29 => x"ef105021",
          30 => x"6f10c061",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef10c065",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"232c4101",
          40 => x"130a0500",
          41 => x"37450000",
          42 => x"1305859b",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"13044100",
          50 => x"ef108063",
          51 => x"37390000",
          52 => x"9309c1ff",
          53 => x"93070400",
          54 => x"13094976",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef100060",
          65 => x"37450000",
          66 => x"1305c59c",
          67 => x"ef10405f",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef10c05c",
          78 => x"37450000",
          79 => x"130545a0",
          80 => x"ef10005c",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74708",
          91 => x"b70600f0",
          92 => x"1377f7fe",
          93 => x"23a2e708",
          94 => x"83a74600",
          95 => x"93c71700",
          96 => x"23a2f600",
          97 => x"67800000",
          98 => x"370700f0",
          99 => x"83274700",
         100 => x"93e70720",
         101 => x"2322f700",
         102 => x"6f000000",
         103 => x"b70700f0",
         104 => x"b70500f0",
         105 => x"370500f0",
         106 => x"9387470f",
         107 => x"9385050f",
         108 => x"83a60700",
         109 => x"03a60500",
         110 => x"03a70700",
         111 => x"e31ad7fe",
         112 => x"b7870100",
         113 => x"b70500f0",
         114 => x"1308f0ff",
         115 => x"9387076a",
         116 => x"23ae050f",
         117 => x"b307f600",
         118 => x"b70600f0",
         119 => x"23ac060f",
         120 => x"33b6c700",
         121 => x"23acf60e",
         122 => x"3306e600",
         123 => x"23aec50e",
         124 => x"83274500",
         125 => x"93c72700",
         126 => x"2322f500",
         127 => x"67800000",
         128 => x"b70700f0",
         129 => x"03a74702",
         130 => x"b70600f0",
         131 => x"93870702",
         132 => x"13774700",
         133 => x"630a0700",
         134 => x"03a74600",
         135 => x"13478700",
         136 => x"23a2e600",
         137 => x"83a78700",
         138 => x"67800000",
         139 => x"b70700f0",
         140 => x"03a7470a",
         141 => x"b70600f0",
         142 => x"1377f7f0",
         143 => x"23a2e70a",
         144 => x"83a74600",
         145 => x"93c74700",
         146 => x"23a2f600",
         147 => x"67800000",
         148 => x"b70700f0",
         149 => x"03a74706",
         150 => x"b70600f0",
         151 => x"137777ff",
         152 => x"23a2e706",
         153 => x"83a74600",
         154 => x"93c70701",
         155 => x"23a2f600",
         156 => x"67800000",
         157 => x"b70700f0",
         158 => x"03a74704",
         159 => x"b70600f0",
         160 => x"137777ff",
         161 => x"23a2e704",
         162 => x"83a74600",
         163 => x"93c70702",
         164 => x"23a2f600",
         165 => x"67800000",
         166 => x"b70700f0",
         167 => x"23ae0700",
         168 => x"03a74700",
         169 => x"13470704",
         170 => x"23a2e700",
         171 => x"67800000",
         172 => x"6f000000",
         173 => x"13050000",
         174 => x"67800000",
         175 => x"13050000",
         176 => x"67800000",
         177 => x"130101f7",
         178 => x"23221100",
         179 => x"23242100",
         180 => x"23263100",
         181 => x"23284100",
         182 => x"232a5100",
         183 => x"232c6100",
         184 => x"232e7100",
         185 => x"23208102",
         186 => x"23229102",
         187 => x"2324a102",
         188 => x"2326b102",
         189 => x"2328c102",
         190 => x"232ad102",
         191 => x"232ce102",
         192 => x"232ef102",
         193 => x"23200105",
         194 => x"23221105",
         195 => x"23242105",
         196 => x"23263105",
         197 => x"23284105",
         198 => x"232a5105",
         199 => x"232c6105",
         200 => x"232e7105",
         201 => x"23208107",
         202 => x"23229107",
         203 => x"2324a107",
         204 => x"2326b107",
         205 => x"2328c107",
         206 => x"232ad107",
         207 => x"232ce107",
         208 => x"232ef107",
         209 => x"f3222034",
         210 => x"23205108",
         211 => x"f3221034",
         212 => x"23225108",
         213 => x"83a20200",
         214 => x"23245108",
         215 => x"f3223034",
         216 => x"23265108",
         217 => x"f3272034",
         218 => x"1307b000",
         219 => x"6374f70c",
         220 => x"37070080",
         221 => x"130797ff",
         222 => x"b387e700",
         223 => x"1307e000",
         224 => x"636ef700",
         225 => x"37370000",
         226 => x"93972700",
         227 => x"13078777",
         228 => x"b387e700",
         229 => x"83a70700",
         230 => x"67800700",
         231 => x"03258102",
         232 => x"83220108",
         233 => x"63c80200",
         234 => x"f3221034",
         235 => x"93824200",
         236 => x"73901234",
         237 => x"832fc107",
         238 => x"032f8107",
         239 => x"832e4107",
         240 => x"032e0107",
         241 => x"832dc106",
         242 => x"032d8106",
         243 => x"832c4106",
         244 => x"032c0106",
         245 => x"832bc105",
         246 => x"032b8105",
         247 => x"832a4105",
         248 => x"032a0105",
         249 => x"8329c104",
         250 => x"03298104",
         251 => x"83284104",
         252 => x"03280104",
         253 => x"8327c103",
         254 => x"03278103",
         255 => x"83264103",
         256 => x"03260103",
         257 => x"8325c102",
         258 => x"83244102",
         259 => x"03240102",
         260 => x"8323c101",
         261 => x"03238101",
         262 => x"83224101",
         263 => x"03220101",
         264 => x"8321c100",
         265 => x"03218100",
         266 => x"83204100",
         267 => x"13010109",
         268 => x"73002030",
         269 => x"93061000",
         270 => x"e3f2f6f6",
         271 => x"e360f7f6",
         272 => x"37370000",
         273 => x"93972700",
         274 => x"1307477b",
         275 => x"b387e700",
         276 => x"83a70700",
         277 => x"67800700",
         278 => x"eff09fdf",
         279 => x"03258102",
         280 => x"6ff01ff4",
         281 => x"eff09fd3",
         282 => x"03258102",
         283 => x"6ff05ff3",
         284 => x"eff09fe2",
         285 => x"03258102",
         286 => x"6ff09ff2",
         287 => x"eff09fce",
         288 => x"03258102",
         289 => x"6ff0dff1",
         290 => x"eff09fd7",
         291 => x"03258102",
         292 => x"6ff01ff1",
         293 => x"eff09fd9",
         294 => x"03258102",
         295 => x"6ff05ff0",
         296 => x"eff05fdd",
         297 => x"03258102",
         298 => x"6ff09fef",
         299 => x"13050100",
         300 => x"eff09fbe",
         301 => x"03258102",
         302 => x"6ff09fee",
         303 => x"9307900a",
         304 => x"6380f814",
         305 => x"63d81703",
         306 => x"9307600d",
         307 => x"638ef818",
         308 => x"938808c0",
         309 => x"9307f000",
         310 => x"63e01705",
         311 => x"b7370000",
         312 => x"9387477e",
         313 => x"93982800",
         314 => x"b388f800",
         315 => x"83a70800",
         316 => x"67800700",
         317 => x"938878fc",
         318 => x"93074002",
         319 => x"63ee1701",
         320 => x"b7470000",
         321 => x"93874782",
         322 => x"93982800",
         323 => x"b388f800",
         324 => x"83a70800",
         325 => x"67800700",
         326 => x"ef10905b",
         327 => x"93078005",
         328 => x"2320f500",
         329 => x"9307f0ff",
         330 => x"13850700",
         331 => x"6ff05fe7",
         332 => x"b7270000",
         333 => x"23a2f500",
         334 => x"93070000",
         335 => x"13850700",
         336 => x"6ff01fe6",
         337 => x"93070000",
         338 => x"13850700",
         339 => x"6ff05fe5",
         340 => x"ef101058",
         341 => x"93079000",
         342 => x"2320f500",
         343 => x"9307f0ff",
         344 => x"13850700",
         345 => x"6ff0dfe3",
         346 => x"ef109056",
         347 => x"9307f001",
         348 => x"2320f500",
         349 => x"9307f0ff",
         350 => x"13850700",
         351 => x"6ff05fe2",
         352 => x"ef101055",
         353 => x"9307d000",
         354 => x"2320f500",
         355 => x"9307f0ff",
         356 => x"13850700",
         357 => x"6ff0dfe0",
         358 => x"ef109053",
         359 => x"93072000",
         360 => x"2320f500",
         361 => x"9307f0ff",
         362 => x"13850700",
         363 => x"6ff05fdf",
         364 => x"13090600",
         365 => x"13840500",
         366 => x"635cc000",
         367 => x"b384c500",
         368 => x"eff09fab",
         369 => x"2300a400",
         370 => x"13041400",
         371 => x"e39a84fe",
         372 => x"13050900",
         373 => x"6ff0dfdc",
         374 => x"13090600",
         375 => x"13840500",
         376 => x"e358c0fe",
         377 => x"b384c500",
         378 => x"03450400",
         379 => x"13041400",
         380 => x"eff0dfa8",
         381 => x"e39a84fe",
         382 => x"13050900",
         383 => x"6ff05fda",
         384 => x"13090000",
         385 => x"93040500",
         386 => x"13040900",
         387 => x"93090900",
         388 => x"93070900",
         389 => x"732410c8",
         390 => x"f32910c0",
         391 => x"f32710c8",
         392 => x"e31af4fe",
         393 => x"37460f00",
         394 => x"13060624",
         395 => x"93060000",
         396 => x"13850900",
         397 => x"93050400",
         398 => x"ef005011",
         399 => x"37460f00",
         400 => x"23a4a400",
         401 => x"13060624",
         402 => x"93060000",
         403 => x"13850900",
         404 => x"93050400",
         405 => x"ef00804c",
         406 => x"23a0a400",
         407 => x"23a2b400",
         408 => x"13050900",
         409 => x"6ff0dfd3",
         410 => x"63180500",
         411 => x"1385819c",
         412 => x"13050500",
         413 => x"6ff0dfd2",
         414 => x"b7870020",
         415 => x"93870700",
         416 => x"13070040",
         417 => x"b387e740",
         418 => x"e364f5fe",
         419 => x"ef105044",
         420 => x"9307c000",
         421 => x"2320f500",
         422 => x"1305f0ff",
         423 => x"13050500",
         424 => x"6ff01fd0",
         425 => x"13030500",
         426 => x"138e0500",
         427 => x"93080000",
         428 => x"63dc0500",
         429 => x"b337a000",
         430 => x"330eb040",
         431 => x"330efe40",
         432 => x"3303a040",
         433 => x"9308f0ff",
         434 => x"63dc0600",
         435 => x"b337c000",
         436 => x"b306d040",
         437 => x"93c8f8ff",
         438 => x"b386f640",
         439 => x"3306c040",
         440 => x"13070600",
         441 => x"13080300",
         442 => x"93070e00",
         443 => x"639c0628",
         444 => x"b7450000",
         445 => x"9385858b",
         446 => x"6376ce0e",
         447 => x"b7060100",
         448 => x"6378d60c",
         449 => x"93360610",
         450 => x"93b61600",
         451 => x"93963600",
         452 => x"3355d600",
         453 => x"b385a500",
         454 => x"83c50500",
         455 => x"13050002",
         456 => x"b386d500",
         457 => x"b305d540",
         458 => x"630cd500",
         459 => x"b317be00",
         460 => x"b356d300",
         461 => x"3317b600",
         462 => x"b3e7f600",
         463 => x"3318b300",
         464 => x"93550701",
         465 => x"33deb702",
         466 => x"13160701",
         467 => x"13560601",
         468 => x"b3f7b702",
         469 => x"13050e00",
         470 => x"3303c603",
         471 => x"93960701",
         472 => x"93570801",
         473 => x"b3e7d700",
         474 => x"63fe6700",
         475 => x"b307f700",
         476 => x"1305feff",
         477 => x"63e8e700",
         478 => x"63f66700",
         479 => x"1305eeff",
         480 => x"b387e700",
         481 => x"b3876740",
         482 => x"33d3b702",
         483 => x"13180801",
         484 => x"13580801",
         485 => x"b3f7b702",
         486 => x"b3066602",
         487 => x"93970701",
         488 => x"3368f800",
         489 => x"93070300",
         490 => x"637cd800",
         491 => x"33080701",
         492 => x"9307f3ff",
         493 => x"6366e800",
         494 => x"6374d800",
         495 => x"9307e3ff",
         496 => x"13150501",
         497 => x"3365f500",
         498 => x"93050000",
         499 => x"6f00000e",
         500 => x"37050001",
         501 => x"93068001",
         502 => x"e37ca6f2",
         503 => x"93060001",
         504 => x"6ff01ff3",
         505 => x"93060000",
         506 => x"630c0600",
         507 => x"b7070100",
         508 => x"637af60c",
         509 => x"93360610",
         510 => x"93b61600",
         511 => x"93963600",
         512 => x"b357d600",
         513 => x"b385f500",
         514 => x"83c70500",
         515 => x"b387d700",
         516 => x"93060002",
         517 => x"b385f640",
         518 => x"6390f60c",
         519 => x"b307ce40",
         520 => x"93051000",
         521 => x"13530701",
         522 => x"b3de6702",
         523 => x"13160701",
         524 => x"13560601",
         525 => x"93560801",
         526 => x"b3f76702",
         527 => x"13850e00",
         528 => x"330ed603",
         529 => x"93970701",
         530 => x"b3e7f600",
         531 => x"63fec701",
         532 => x"b307f700",
         533 => x"1385feff",
         534 => x"63e8e700",
         535 => x"63f6c701",
         536 => x"1385eeff",
         537 => x"b387e700",
         538 => x"b387c741",
         539 => x"33de6702",
         540 => x"13180801",
         541 => x"13580801",
         542 => x"b3f76702",
         543 => x"b306c603",
         544 => x"93970701",
         545 => x"3368f800",
         546 => x"93070e00",
         547 => x"637cd800",
         548 => x"33080701",
         549 => x"9307feff",
         550 => x"6366e800",
         551 => x"6374d800",
         552 => x"9307eeff",
         553 => x"13150501",
         554 => x"3365f500",
         555 => x"638a0800",
         556 => x"b337a000",
         557 => x"b305b040",
         558 => x"b385f540",
         559 => x"3305a040",
         560 => x"67800000",
         561 => x"b7070001",
         562 => x"93068001",
         563 => x"e37af6f2",
         564 => x"93060001",
         565 => x"6ff0dff2",
         566 => x"3317b600",
         567 => x"b356fe00",
         568 => x"13550701",
         569 => x"331ebe00",
         570 => x"b357f300",
         571 => x"b3e7c701",
         572 => x"33dea602",
         573 => x"13160701",
         574 => x"13560601",
         575 => x"3318b300",
         576 => x"b3f6a602",
         577 => x"3303c603",
         578 => x"93950601",
         579 => x"93d60701",
         580 => x"b3e6b600",
         581 => x"93050e00",
         582 => x"63fe6600",
         583 => x"b306d700",
         584 => x"9305feff",
         585 => x"63e8e600",
         586 => x"63f66600",
         587 => x"9305eeff",
         588 => x"b386e600",
         589 => x"b3866640",
         590 => x"33d3a602",
         591 => x"93970701",
         592 => x"93d70701",
         593 => x"b3f6a602",
         594 => x"33066602",
         595 => x"93960601",
         596 => x"b3e7d700",
         597 => x"93060300",
         598 => x"63fec700",
         599 => x"b307f700",
         600 => x"9306f3ff",
         601 => x"63e8e700",
         602 => x"63f6c700",
         603 => x"9306e3ff",
         604 => x"b387e700",
         605 => x"93950501",
         606 => x"b387c740",
         607 => x"b3e5d500",
         608 => x"6ff05fea",
         609 => x"6366de18",
         610 => x"b7070100",
         611 => x"63f4f604",
         612 => x"13b70610",
         613 => x"13371700",
         614 => x"13173700",
         615 => x"b7470000",
         616 => x"b3d5e600",
         617 => x"9387878b",
         618 => x"b387b700",
         619 => x"83c70700",
         620 => x"b387e700",
         621 => x"13070002",
         622 => x"b305f740",
         623 => x"6316f702",
         624 => x"13051000",
         625 => x"e3e4c6ef",
         626 => x"3335c300",
         627 => x"13351500",
         628 => x"6ff0dfed",
         629 => x"b7070001",
         630 => x"13078001",
         631 => x"e3f0f6fc",
         632 => x"13070001",
         633 => x"6ff09ffb",
         634 => x"3357f600",
         635 => x"b396b600",
         636 => x"b366d700",
         637 => x"3357fe00",
         638 => x"331ebe00",
         639 => x"b357f300",
         640 => x"b3e7c701",
         641 => x"13de0601",
         642 => x"335fc703",
         643 => x"13980601",
         644 => x"13580801",
         645 => x"3316b600",
         646 => x"3377c703",
         647 => x"b30ee803",
         648 => x"13150701",
         649 => x"13d70701",
         650 => x"3367a700",
         651 => x"13050f00",
         652 => x"637ed701",
         653 => x"3387e600",
         654 => x"1305ffff",
         655 => x"6368d700",
         656 => x"6376d701",
         657 => x"1305efff",
         658 => x"3307d700",
         659 => x"3307d741",
         660 => x"b35ec703",
         661 => x"93970701",
         662 => x"93d70701",
         663 => x"3377c703",
         664 => x"3308d803",
         665 => x"13170701",
         666 => x"b3e7e700",
         667 => x"13870e00",
         668 => x"63fe0701",
         669 => x"b387f600",
         670 => x"1387feff",
         671 => x"63e8d700",
         672 => x"63f60701",
         673 => x"1387eeff",
         674 => x"b387d700",
         675 => x"13150501",
         676 => x"b70e0100",
         677 => x"3365e500",
         678 => x"9386feff",
         679 => x"3377d500",
         680 => x"b3870741",
         681 => x"b376d600",
         682 => x"13580501",
         683 => x"13560601",
         684 => x"330ed702",
         685 => x"b306d802",
         686 => x"3307c702",
         687 => x"3308c802",
         688 => x"3306d700",
         689 => x"13570e01",
         690 => x"3307c700",
         691 => x"6374d700",
         692 => x"3308d801",
         693 => x"93560701",
         694 => x"b3860601",
         695 => x"63e6d702",
         696 => x"e394d7ce",
         697 => x"b7070100",
         698 => x"9387f7ff",
         699 => x"3377f700",
         700 => x"13170701",
         701 => x"337efe00",
         702 => x"3313b300",
         703 => x"3307c701",
         704 => x"93050000",
         705 => x"e374e3da",
         706 => x"1305f5ff",
         707 => x"6ff0dfcb",
         708 => x"93050000",
         709 => x"13050000",
         710 => x"6ff05fd9",
         711 => x"93080500",
         712 => x"13830500",
         713 => x"13070600",
         714 => x"13080500",
         715 => x"93870500",
         716 => x"63920628",
         717 => x"b7450000",
         718 => x"9385858b",
         719 => x"6376c30e",
         720 => x"b7060100",
         721 => x"6378d60c",
         722 => x"93360610",
         723 => x"93b61600",
         724 => x"93963600",
         725 => x"3355d600",
         726 => x"b385a500",
         727 => x"83c50500",
         728 => x"13050002",
         729 => x"b386d500",
         730 => x"b305d540",
         731 => x"630cd500",
         732 => x"b317b300",
         733 => x"b3d6d800",
         734 => x"3317b600",
         735 => x"b3e7f600",
         736 => x"3398b800",
         737 => x"93550701",
         738 => x"33d3b702",
         739 => x"13160701",
         740 => x"13560601",
         741 => x"b3f7b702",
         742 => x"13050300",
         743 => x"b3086602",
         744 => x"93960701",
         745 => x"93570801",
         746 => x"b3e7d700",
         747 => x"63fe1701",
         748 => x"b307f700",
         749 => x"1305f3ff",
         750 => x"63e8e700",
         751 => x"63f61701",
         752 => x"1305e3ff",
         753 => x"b387e700",
         754 => x"b3871741",
         755 => x"b3d8b702",
         756 => x"13180801",
         757 => x"13580801",
         758 => x"b3f7b702",
         759 => x"b3061603",
         760 => x"93970701",
         761 => x"3368f800",
         762 => x"93870800",
         763 => x"637cd800",
         764 => x"33080701",
         765 => x"9387f8ff",
         766 => x"6366e800",
         767 => x"6374d800",
         768 => x"9387e8ff",
         769 => x"13150501",
         770 => x"3365f500",
         771 => x"93050000",
         772 => x"67800000",
         773 => x"37050001",
         774 => x"93068001",
         775 => x"e37ca6f2",
         776 => x"93060001",
         777 => x"6ff01ff3",
         778 => x"93060000",
         779 => x"630c0600",
         780 => x"b7070100",
         781 => x"6370f60c",
         782 => x"93360610",
         783 => x"93b61600",
         784 => x"93963600",
         785 => x"b357d600",
         786 => x"b385f500",
         787 => x"83c70500",
         788 => x"b387d700",
         789 => x"93060002",
         790 => x"b385f640",
         791 => x"6396f60a",
         792 => x"b307c340",
         793 => x"93051000",
         794 => x"93580701",
         795 => x"33de1703",
         796 => x"13160701",
         797 => x"13560601",
         798 => x"93560801",
         799 => x"b3f71703",
         800 => x"13050e00",
         801 => x"3303c603",
         802 => x"93970701",
         803 => x"b3e7f600",
         804 => x"63fe6700",
         805 => x"b307f700",
         806 => x"1305feff",
         807 => x"63e8e700",
         808 => x"63f66700",
         809 => x"1305eeff",
         810 => x"b387e700",
         811 => x"b3876740",
         812 => x"33d31703",
         813 => x"13180801",
         814 => x"13580801",
         815 => x"b3f71703",
         816 => x"b3066602",
         817 => x"93970701",
         818 => x"3368f800",
         819 => x"93070300",
         820 => x"637cd800",
         821 => x"33080701",
         822 => x"9307f3ff",
         823 => x"6366e800",
         824 => x"6374d800",
         825 => x"9307e3ff",
         826 => x"13150501",
         827 => x"3365f500",
         828 => x"67800000",
         829 => x"b7070001",
         830 => x"93068001",
         831 => x"e374f6f4",
         832 => x"93060001",
         833 => x"6ff01ff4",
         834 => x"3317b600",
         835 => x"b356f300",
         836 => x"13550701",
         837 => x"3313b300",
         838 => x"b3d7f800",
         839 => x"b3e76700",
         840 => x"33d3a602",
         841 => x"13160701",
         842 => x"13560601",
         843 => x"3398b800",
         844 => x"b3f6a602",
         845 => x"b3086602",
         846 => x"93950601",
         847 => x"93d60701",
         848 => x"b3e6b600",
         849 => x"93050300",
         850 => x"63fe1601",
         851 => x"b306d700",
         852 => x"9305f3ff",
         853 => x"63e8e600",
         854 => x"63f61601",
         855 => x"9305e3ff",
         856 => x"b386e600",
         857 => x"b3861641",
         858 => x"b3d8a602",
         859 => x"93970701",
         860 => x"93d70701",
         861 => x"b3f6a602",
         862 => x"33061603",
         863 => x"93960601",
         864 => x"b3e7d700",
         865 => x"93860800",
         866 => x"63fec700",
         867 => x"b307f700",
         868 => x"9386f8ff",
         869 => x"63e8e700",
         870 => x"63f6c700",
         871 => x"9386e8ff",
         872 => x"b387e700",
         873 => x"93950501",
         874 => x"b387c740",
         875 => x"b3e5d500",
         876 => x"6ff09feb",
         877 => x"63e6d518",
         878 => x"b7070100",
         879 => x"63f4f604",
         880 => x"13b70610",
         881 => x"13371700",
         882 => x"13173700",
         883 => x"b7470000",
         884 => x"b3d5e600",
         885 => x"9387878b",
         886 => x"b387b700",
         887 => x"83c70700",
         888 => x"b387e700",
         889 => x"13070002",
         890 => x"b305f740",
         891 => x"6316f702",
         892 => x"13051000",
         893 => x"e3ee66e0",
         894 => x"33b5c800",
         895 => x"13351500",
         896 => x"67800000",
         897 => x"b7070001",
         898 => x"13078001",
         899 => x"e3f0f6fc",
         900 => x"13070001",
         901 => x"6ff09ffb",
         902 => x"3357f600",
         903 => x"b396b600",
         904 => x"b366d700",
         905 => x"3357f300",
         906 => x"3313b300",
         907 => x"b3d7f800",
         908 => x"b3e76700",
         909 => x"13d30601",
         910 => x"b35e6702",
         911 => x"13980601",
         912 => x"13580801",
         913 => x"3316b600",
         914 => x"33776702",
         915 => x"330ed803",
         916 => x"13150701",
         917 => x"13d70701",
         918 => x"3367a700",
         919 => x"13850e00",
         920 => x"637ec701",
         921 => x"3387e600",
         922 => x"1385feff",
         923 => x"6368d700",
         924 => x"6376c701",
         925 => x"1385eeff",
         926 => x"3307d700",
         927 => x"3307c741",
         928 => x"335e6702",
         929 => x"93970701",
         930 => x"93d70701",
         931 => x"33776702",
         932 => x"3308c803",
         933 => x"13170701",
         934 => x"b3e7e700",
         935 => x"13070e00",
         936 => x"63fe0701",
         937 => x"b387f600",
         938 => x"1307feff",
         939 => x"63e8d700",
         940 => x"63f60701",
         941 => x"1307eeff",
         942 => x"b387d700",
         943 => x"13150501",
         944 => x"370e0100",
         945 => x"3365e500",
         946 => x"9306feff",
         947 => x"3377d500",
         948 => x"b3870741",
         949 => x"b376d600",
         950 => x"13580501",
         951 => x"13560601",
         952 => x"3303d702",
         953 => x"b306d802",
         954 => x"3307c702",
         955 => x"3308c802",
         956 => x"3306d700",
         957 => x"13570301",
         958 => x"3307c700",
         959 => x"6374d700",
         960 => x"3308c801",
         961 => x"93560701",
         962 => x"b3860601",
         963 => x"63e6d702",
         964 => x"e39ed7ce",
         965 => x"b7070100",
         966 => x"9387f7ff",
         967 => x"3377f700",
         968 => x"13170701",
         969 => x"3373f300",
         970 => x"b398b800",
         971 => x"33076700",
         972 => x"93050000",
         973 => x"e3fee8cc",
         974 => x"1305f5ff",
         975 => x"6ff01fcd",
         976 => x"93050000",
         977 => x"13050000",
         978 => x"67800000",
         979 => x"13080600",
         980 => x"93070500",
         981 => x"13870500",
         982 => x"63960620",
         983 => x"b7480000",
         984 => x"9388888b",
         985 => x"63fcc50c",
         986 => x"b7060100",
         987 => x"637ed60a",
         988 => x"93360610",
         989 => x"93b61600",
         990 => x"93963600",
         991 => x"3353d600",
         992 => x"b3886800",
         993 => x"83c80800",
         994 => x"13030002",
         995 => x"b386d800",
         996 => x"b308d340",
         997 => x"630cd300",
         998 => x"33971501",
         999 => x"b356d500",
        1000 => x"33181601",
        1001 => x"33e7e600",
        1002 => x"b3171501",
        1003 => x"13560801",
        1004 => x"b356c702",
        1005 => x"13150801",
        1006 => x"13550501",
        1007 => x"3377c702",
        1008 => x"b386a602",
        1009 => x"93150701",
        1010 => x"13d70701",
        1011 => x"3367b700",
        1012 => x"637ad700",
        1013 => x"3307e800",
        1014 => x"63660701",
        1015 => x"6374d700",
        1016 => x"33070701",
        1017 => x"3307d740",
        1018 => x"b356c702",
        1019 => x"3377c702",
        1020 => x"b386a602",
        1021 => x"93970701",
        1022 => x"13170701",
        1023 => x"93d70701",
        1024 => x"b3e7e700",
        1025 => x"63fad700",
        1026 => x"b307f800",
        1027 => x"63e60701",
        1028 => x"63f4d700",
        1029 => x"b3870701",
        1030 => x"b387d740",
        1031 => x"33d51701",
        1032 => x"93050000",
        1033 => x"67800000",
        1034 => x"37030001",
        1035 => x"93068001",
        1036 => x"e37666f4",
        1037 => x"93060001",
        1038 => x"6ff05ff4",
        1039 => x"93060000",
        1040 => x"630c0600",
        1041 => x"37070100",
        1042 => x"637ee606",
        1043 => x"93360610",
        1044 => x"93b61600",
        1045 => x"93963600",
        1046 => x"3357d600",
        1047 => x"b388e800",
        1048 => x"03c70800",
        1049 => x"3307d700",
        1050 => x"93060002",
        1051 => x"b388e640",
        1052 => x"6394e606",
        1053 => x"3387c540",
        1054 => x"93550801",
        1055 => x"3356b702",
        1056 => x"13150801",
        1057 => x"13550501",
        1058 => x"93d60701",
        1059 => x"3377b702",
        1060 => x"3306a602",
        1061 => x"13170701",
        1062 => x"33e7e600",
        1063 => x"637ac700",
        1064 => x"3307e800",
        1065 => x"63660701",
        1066 => x"6374c700",
        1067 => x"33070701",
        1068 => x"3307c740",
        1069 => x"b356b702",
        1070 => x"3377b702",
        1071 => x"b386a602",
        1072 => x"6ff05ff3",
        1073 => x"37070001",
        1074 => x"93068001",
        1075 => x"e376e6f8",
        1076 => x"93060001",
        1077 => x"6ff05ff8",
        1078 => x"33181601",
        1079 => x"b3d6e500",
        1080 => x"b3171501",
        1081 => x"b3951501",
        1082 => x"3357e500",
        1083 => x"13550801",
        1084 => x"3367b700",
        1085 => x"b3d5a602",
        1086 => x"13130801",
        1087 => x"13530301",
        1088 => x"b3f6a602",
        1089 => x"b3856502",
        1090 => x"13960601",
        1091 => x"93560701",
        1092 => x"b3e6c600",
        1093 => x"63fab600",
        1094 => x"b306d800",
        1095 => x"63e60601",
        1096 => x"63f4b600",
        1097 => x"b3860601",
        1098 => x"b386b640",
        1099 => x"33d6a602",
        1100 => x"13170701",
        1101 => x"13570701",
        1102 => x"b3f6a602",
        1103 => x"33066602",
        1104 => x"93960601",
        1105 => x"3367d700",
        1106 => x"637ac700",
        1107 => x"3307e800",
        1108 => x"63660701",
        1109 => x"6374c700",
        1110 => x"33070701",
        1111 => x"3307c740",
        1112 => x"6ff09ff1",
        1113 => x"63e4d51c",
        1114 => x"37080100",
        1115 => x"63fe0605",
        1116 => x"13b80610",
        1117 => x"13381800",
        1118 => x"13183800",
        1119 => x"b7480000",
        1120 => x"33d30601",
        1121 => x"9388888b",
        1122 => x"b3886800",
        1123 => x"83c80800",
        1124 => x"13030002",
        1125 => x"b3880801",
        1126 => x"33081341",
        1127 => x"63101305",
        1128 => x"63e4b600",
        1129 => x"636cc500",
        1130 => x"3306c540",
        1131 => x"b386d540",
        1132 => x"3337c500",
        1133 => x"93070600",
        1134 => x"3387e640",
        1135 => x"13850700",
        1136 => x"93050700",
        1137 => x"67800000",
        1138 => x"b7080001",
        1139 => x"13088001",
        1140 => x"e3f616fb",
        1141 => x"13080001",
        1142 => x"6ff05ffa",
        1143 => x"b3571601",
        1144 => x"b3960601",
        1145 => x"b3e6d700",
        1146 => x"33d71501",
        1147 => x"13de0601",
        1148 => x"335fc703",
        1149 => x"13930601",
        1150 => x"13530301",
        1151 => x"b3970501",
        1152 => x"b3551501",
        1153 => x"b3e5f500",
        1154 => x"93d70501",
        1155 => x"33160601",
        1156 => x"33150501",
        1157 => x"3377c703",
        1158 => x"b30ee303",
        1159 => x"13170701",
        1160 => x"b3e7e700",
        1161 => x"13070f00",
        1162 => x"63fed701",
        1163 => x"b387f600",
        1164 => x"1307ffff",
        1165 => x"63e8d700",
        1166 => x"63f6d701",
        1167 => x"1307efff",
        1168 => x"b387d700",
        1169 => x"b387d741",
        1170 => x"b3dec703",
        1171 => x"93950501",
        1172 => x"93d50501",
        1173 => x"b3f7c703",
        1174 => x"138e0e00",
        1175 => x"3303d303",
        1176 => x"93970701",
        1177 => x"b3e5f500",
        1178 => x"63fe6500",
        1179 => x"b385b600",
        1180 => x"138efeff",
        1181 => x"63e8d500",
        1182 => x"63f66500",
        1183 => x"138eeeff",
        1184 => x"b385d500",
        1185 => x"93170701",
        1186 => x"370f0100",
        1187 => x"b3e7c701",
        1188 => x"b3856540",
        1189 => x"1303ffff",
        1190 => x"33f76700",
        1191 => x"135e0601",
        1192 => x"93d70701",
        1193 => x"33736600",
        1194 => x"b30e6702",
        1195 => x"33836702",
        1196 => x"3307c703",
        1197 => x"b387c703",
        1198 => x"330e6700",
        1199 => x"13d70e01",
        1200 => x"3307c701",
        1201 => x"63746700",
        1202 => x"b387e701",
        1203 => x"13530701",
        1204 => x"b307f300",
        1205 => x"37030100",
        1206 => x"1303f3ff",
        1207 => x"33776700",
        1208 => x"13170701",
        1209 => x"b3fe6e00",
        1210 => x"3307d701",
        1211 => x"63e6f500",
        1212 => x"639ef500",
        1213 => x"637ce500",
        1214 => x"3306c740",
        1215 => x"3333c700",
        1216 => x"b306d300",
        1217 => x"13070600",
        1218 => x"b387d740",
        1219 => x"3307e540",
        1220 => x"3335e500",
        1221 => x"b385f540",
        1222 => x"b385a540",
        1223 => x"b3981501",
        1224 => x"33570701",
        1225 => x"33e5e800",
        1226 => x"b3d50501",
        1227 => x"67800000",
        1228 => x"13030500",
        1229 => x"630a0600",
        1230 => x"2300b300",
        1231 => x"1306f6ff",
        1232 => x"13031300",
        1233 => x"e31a06fe",
        1234 => x"67800000",
        1235 => x"13030500",
        1236 => x"630e0600",
        1237 => x"83830500",
        1238 => x"23007300",
        1239 => x"1306f6ff",
        1240 => x"13031300",
        1241 => x"93851500",
        1242 => x"e31606fe",
        1243 => x"67800000",
        1244 => x"630c0602",
        1245 => x"13030500",
        1246 => x"93061000",
        1247 => x"636ab500",
        1248 => x"9306f0ff",
        1249 => x"1307f6ff",
        1250 => x"3303e300",
        1251 => x"b385e500",
        1252 => x"83830500",
        1253 => x"23007300",
        1254 => x"1306f6ff",
        1255 => x"3303d300",
        1256 => x"b385d500",
        1257 => x"e31606fe",
        1258 => x"67800000",
        1259 => x"6f000000",
        1260 => x"130101ff",
        1261 => x"23248100",
        1262 => x"13040000",
        1263 => x"23229100",
        1264 => x"23202101",
        1265 => x"23261100",
        1266 => x"93040500",
        1267 => x"13090400",
        1268 => x"93070400",
        1269 => x"732410c8",
        1270 => x"732910c0",
        1271 => x"f32710c8",
        1272 => x"e31af4fe",
        1273 => x"37460f00",
        1274 => x"13060624",
        1275 => x"93060000",
        1276 => x"13050900",
        1277 => x"93050400",
        1278 => x"eff05fb5",
        1279 => x"37460f00",
        1280 => x"23a4a400",
        1281 => x"93050400",
        1282 => x"13050900",
        1283 => x"13060624",
        1284 => x"93060000",
        1285 => x"eff08ff0",
        1286 => x"8320c100",
        1287 => x"03248100",
        1288 => x"23a0a400",
        1289 => x"23a2b400",
        1290 => x"03290100",
        1291 => x"83244100",
        1292 => x"13050000",
        1293 => x"13010101",
        1294 => x"67800000",
        1295 => x"13050000",
        1296 => x"67800000",
        1297 => x"13050000",
        1298 => x"67800000",
        1299 => x"130101ff",
        1300 => x"23202101",
        1301 => x"23261100",
        1302 => x"13090600",
        1303 => x"6356c002",
        1304 => x"23248100",
        1305 => x"23229100",
        1306 => x"13840500",
        1307 => x"b384c500",
        1308 => x"03450400",
        1309 => x"13041400",
        1310 => x"efe05fc0",
        1311 => x"e39a84fe",
        1312 => x"03248100",
        1313 => x"83244100",
        1314 => x"8320c100",
        1315 => x"13050900",
        1316 => x"03290100",
        1317 => x"13010101",
        1318 => x"67800000",
        1319 => x"130101ff",
        1320 => x"23202101",
        1321 => x"23261100",
        1322 => x"13090600",
        1323 => x"6356c002",
        1324 => x"23248100",
        1325 => x"23229100",
        1326 => x"13840500",
        1327 => x"b384c500",
        1328 => x"efe09fbb",
        1329 => x"13041400",
        1330 => x"a30fa4fe",
        1331 => x"e39a84fe",
        1332 => x"03248100",
        1333 => x"83244100",
        1334 => x"8320c100",
        1335 => x"13050900",
        1336 => x"03290100",
        1337 => x"13010101",
        1338 => x"67800000",
        1339 => x"13051000",
        1340 => x"67800000",
        1341 => x"130101ff",
        1342 => x"23261100",
        1343 => x"ef00505d",
        1344 => x"8320c100",
        1345 => x"93076001",
        1346 => x"2320f500",
        1347 => x"1305f0ff",
        1348 => x"13010101",
        1349 => x"67800000",
        1350 => x"1305f0ff",
        1351 => x"67800000",
        1352 => x"b7270000",
        1353 => x"23a2f500",
        1354 => x"13050000",
        1355 => x"67800000",
        1356 => x"13051000",
        1357 => x"67800000",
        1358 => x"13050000",
        1359 => x"67800000",
        1360 => x"130101fe",
        1361 => x"2324c100",
        1362 => x"2326d100",
        1363 => x"2328e100",
        1364 => x"232af100",
        1365 => x"232c0101",
        1366 => x"232e1101",
        1367 => x"1305f0ff",
        1368 => x"13010102",
        1369 => x"67800000",
        1370 => x"130101ff",
        1371 => x"23261100",
        1372 => x"ef001056",
        1373 => x"8320c100",
        1374 => x"9307a000",
        1375 => x"2320f500",
        1376 => x"1305f0ff",
        1377 => x"13010101",
        1378 => x"67800000",
        1379 => x"130101ff",
        1380 => x"23261100",
        1381 => x"ef00d053",
        1382 => x"8320c100",
        1383 => x"93072000",
        1384 => x"2320f500",
        1385 => x"1305f0ff",
        1386 => x"13010101",
        1387 => x"67800000",
        1388 => x"b7270000",
        1389 => x"23a2f500",
        1390 => x"13050000",
        1391 => x"67800000",
        1392 => x"130101ff",
        1393 => x"23261100",
        1394 => x"ef009050",
        1395 => x"8320c100",
        1396 => x"9307f001",
        1397 => x"2320f500",
        1398 => x"1305f0ff",
        1399 => x"13010101",
        1400 => x"67800000",
        1401 => x"130101ff",
        1402 => x"23261100",
        1403 => x"ef00504e",
        1404 => x"8320c100",
        1405 => x"9307b000",
        1406 => x"2320f500",
        1407 => x"1305f0ff",
        1408 => x"13010101",
        1409 => x"67800000",
        1410 => x"130101ff",
        1411 => x"23261100",
        1412 => x"ef00104c",
        1413 => x"8320c100",
        1414 => x"9307c000",
        1415 => x"2320f500",
        1416 => x"1305f0ff",
        1417 => x"13010101",
        1418 => x"67800000",
        1419 => x"03a7c187",
        1420 => x"b7870020",
        1421 => x"93870700",
        1422 => x"93060040",
        1423 => x"b387d740",
        1424 => x"630c0700",
        1425 => x"3305a700",
        1426 => x"63e2a702",
        1427 => x"23aea186",
        1428 => x"13050700",
        1429 => x"67800000",
        1430 => x"9386819c",
        1431 => x"1387819c",
        1432 => x"23aed186",
        1433 => x"3305a700",
        1434 => x"e3f2a7fe",
        1435 => x"130101ff",
        1436 => x"23261100",
        1437 => x"ef00d045",
        1438 => x"8320c100",
        1439 => x"9307c000",
        1440 => x"2320f500",
        1441 => x"1307f0ff",
        1442 => x"13050700",
        1443 => x"13010101",
        1444 => x"67800000",
        1445 => x"370700f0",
        1446 => x"13070702",
        1447 => x"83274700",
        1448 => x"93f74700",
        1449 => x"e38c07fe",
        1450 => x"03258700",
        1451 => x"1375f50f",
        1452 => x"67800000",
        1453 => x"f32710fc",
        1454 => x"63960700",
        1455 => x"b7f7fa02",
        1456 => x"93870708",
        1457 => x"63060500",
        1458 => x"33d5a702",
        1459 => x"1305f5ff",
        1460 => x"b70700f0",
        1461 => x"23a6a702",
        1462 => x"23a0b702",
        1463 => x"67800000",
        1464 => x"370700f0",
        1465 => x"1375f50f",
        1466 => x"13070702",
        1467 => x"2324a700",
        1468 => x"83274700",
        1469 => x"93f70701",
        1470 => x"e38c07fe",
        1471 => x"67800000",
        1472 => x"630e0502",
        1473 => x"130101ff",
        1474 => x"23248100",
        1475 => x"23261100",
        1476 => x"13040500",
        1477 => x"03450500",
        1478 => x"630a0500",
        1479 => x"13041400",
        1480 => x"eff01ffc",
        1481 => x"03450400",
        1482 => x"e31a05fe",
        1483 => x"8320c100",
        1484 => x"03248100",
        1485 => x"13010101",
        1486 => x"67800000",
        1487 => x"67800000",
        1488 => x"130101f9",
        1489 => x"23248106",
        1490 => x"23229106",
        1491 => x"23261106",
        1492 => x"23202107",
        1493 => x"232e3105",
        1494 => x"232c4105",
        1495 => x"232a5105",
        1496 => x"23286105",
        1497 => x"23267105",
        1498 => x"23248105",
        1499 => x"23229105",
        1500 => x"2320a105",
        1501 => x"93040500",
        1502 => x"13840500",
        1503 => x"232c0100",
        1504 => x"232e0100",
        1505 => x"23200102",
        1506 => x"23220102",
        1507 => x"23240102",
        1508 => x"23260102",
        1509 => x"23280102",
        1510 => x"232a0102",
        1511 => x"232c0102",
        1512 => x"232e0102",
        1513 => x"97f2ffff",
        1514 => x"938202b2",
        1515 => x"73905230",
        1516 => x"37c50100",
        1517 => x"93050004",
        1518 => x"13050520",
        1519 => x"eff09fef",
        1520 => x"f32710fc",
        1521 => x"93d71700",
        1522 => x"370700f0",
        1523 => x"9387f7ff",
        1524 => x"2326f708",
        1525 => x"93051001",
        1526 => x"2320b708",
        1527 => x"732710fc",
        1528 => x"b7270000",
        1529 => x"93870771",
        1530 => x"3357f702",
        1531 => x"37260000",
        1532 => x"b70700f0",
        1533 => x"1306f670",
        1534 => x"b70600f0",
        1535 => x"1307f7ff",
        1536 => x"23a8e70a",
        1537 => x"23a6c70a",
        1538 => x"23a0b70a",
        1539 => x"93078070",
        1540 => x"23a0f606",
        1541 => x"f32710fc",
        1542 => x"37571200",
        1543 => x"130707f8",
        1544 => x"b3d7e702",
        1545 => x"370700f0",
        1546 => x"9387f7ff",
        1547 => x"93970701",
        1548 => x"93e78700",
        1549 => x"2320f704",
        1550 => x"b70700f0",
        1551 => x"1307a007",
        1552 => x"23ace700",
        1553 => x"93020008",
        1554 => x"73904230",
        1555 => x"b7220000",
        1556 => x"93828280",
        1557 => x"73900230",
        1558 => x"b7490000",
        1559 => x"138549a0",
        1560 => x"eff01fea",
        1561 => x"63549002",
        1562 => x"1389f4ff",
        1563 => x"9304f0ff",
        1564 => x"03250400",
        1565 => x"1309f9ff",
        1566 => x"13044400",
        1567 => x"eff05fe8",
        1568 => x"138549a0",
        1569 => x"eff0dfe7",
        1570 => x"e31499fe",
        1571 => x"37450000",
        1572 => x"1305859d",
        1573 => x"37f9eeee",
        1574 => x"b7faeeee",
        1575 => x"b7090010",
        1576 => x"37140000",
        1577 => x"eff0dfe5",
        1578 => x"374b0000",
        1579 => x"9389f9ff",
        1580 => x"1309f9ee",
        1581 => x"938aeaee",
        1582 => x"130404e1",
        1583 => x"93040000",
        1584 => x"b71b0000",
        1585 => x"938b0b2c",
        1586 => x"130af000",
        1587 => x"6f00c000",
        1588 => x"938bfbff",
        1589 => x"63840b18",
        1590 => x"93050000",
        1591 => x"13058100",
        1592 => x"ef005029",
        1593 => x"e31605fe",
        1594 => x"032c8100",
        1595 => x"8325c100",
        1596 => x"13060400",
        1597 => x"9357cc01",
        1598 => x"13974500",
        1599 => x"b367f700",
        1600 => x"b3f73701",
        1601 => x"33773c01",
        1602 => x"13d5f541",
        1603 => x"13d88501",
        1604 => x"3307f700",
        1605 => x"33070701",
        1606 => x"9377d500",
        1607 => x"3307f700",
        1608 => x"33774703",
        1609 => x"937725ff",
        1610 => x"93860400",
        1611 => x"13050c00",
        1612 => x"938bfbff",
        1613 => x"3307f700",
        1614 => x"b307ec40",
        1615 => x"1357f741",
        1616 => x"3338fc00",
        1617 => x"3387e540",
        1618 => x"33070741",
        1619 => x"b3885703",
        1620 => x"33072703",
        1621 => x"33b82703",
        1622 => x"33071701",
        1623 => x"b3872703",
        1624 => x"33070701",
        1625 => x"1358f741",
        1626 => x"13783800",
        1627 => x"b307f800",
        1628 => x"33b80701",
        1629 => x"3307e800",
        1630 => x"1318e701",
        1631 => x"93d72700",
        1632 => x"b367f800",
        1633 => x"13582740",
        1634 => x"93184800",
        1635 => x"13d3c701",
        1636 => x"33e36800",
        1637 => x"33733301",
        1638 => x"b3f83701",
        1639 => x"135e8801",
        1640 => x"1357f741",
        1641 => x"b3886800",
        1642 => x"b388c801",
        1643 => x"1373d700",
        1644 => x"b3886800",
        1645 => x"b3f84803",
        1646 => x"137727ff",
        1647 => x"939c4700",
        1648 => x"b38cfc40",
        1649 => x"939c2c00",
        1650 => x"b30c9c41",
        1651 => x"b388e800",
        1652 => x"33871741",
        1653 => x"93d8f841",
        1654 => x"33b3e700",
        1655 => x"33081841",
        1656 => x"33086840",
        1657 => x"33082803",
        1658 => x"33035703",
        1659 => x"b3382703",
        1660 => x"33086800",
        1661 => x"33072703",
        1662 => x"33081801",
        1663 => x"9358f841",
        1664 => x"93f83800",
        1665 => x"3387e800",
        1666 => x"b3381701",
        1667 => x"b3880801",
        1668 => x"9398e801",
        1669 => x"13572700",
        1670 => x"33e7e800",
        1671 => x"13184700",
        1672 => x"3307e840",
        1673 => x"13172700",
        1674 => x"338de740",
        1675 => x"efe09fc7",
        1676 => x"83260101",
        1677 => x"13070500",
        1678 => x"13880c00",
        1679 => x"93070d00",
        1680 => x"13060c00",
        1681 => x"93058ba0",
        1682 => x"13058101",
        1683 => x"ef008044",
        1684 => x"13058101",
        1685 => x"eff0dfca",
        1686 => x"e3900be8",
        1687 => x"73001000",
        1688 => x"370700f0",
        1689 => x"9306f00f",
        1690 => x"b70700f0",
        1691 => x"2324d706",
        1692 => x"03a70704",
        1693 => x"13670730",
        1694 => x"23a0e704",
        1695 => x"13070009",
        1696 => x"23a4e704",
        1697 => x"6ff0dfe3",
        1698 => x"130101ff",
        1699 => x"23248100",
        1700 => x"23261100",
        1701 => x"93070000",
        1702 => x"13040500",
        1703 => x"63880700",
        1704 => x"93050000",
        1705 => x"97000000",
        1706 => x"e7000000",
        1707 => x"83a70188",
        1708 => x"63840700",
        1709 => x"e7800700",
        1710 => x"13050400",
        1711 => x"eff01f8f",
        1712 => x"13050000",
        1713 => x"67800000",
        1714 => x"130101ff",
        1715 => x"23248100",
        1716 => x"23261100",
        1717 => x"13040500",
        1718 => x"2316b500",
        1719 => x"2317c500",
        1720 => x"23200500",
        1721 => x"23220500",
        1722 => x"23240500",
        1723 => x"23220506",
        1724 => x"23280500",
        1725 => x"232a0500",
        1726 => x"232c0500",
        1727 => x"13068000",
        1728 => x"93050000",
        1729 => x"1305c505",
        1730 => x"eff09f82",
        1731 => x"b7270000",
        1732 => x"938747f0",
        1733 => x"2322f402",
        1734 => x"b7270000",
        1735 => x"9387c7f5",
        1736 => x"2324f402",
        1737 => x"b7270000",
        1738 => x"938707fe",
        1739 => x"2326f402",
        1740 => x"b7270000",
        1741 => x"93878703",
        1742 => x"8320c100",
        1743 => x"23208402",
        1744 => x"2328f402",
        1745 => x"03248100",
        1746 => x"13010101",
        1747 => x"67800000",
        1748 => x"b7350000",
        1749 => x"37050020",
        1750 => x"13868181",
        1751 => x"9385054b",
        1752 => x"13054502",
        1753 => x"6f00c021",
        1754 => x"83254500",
        1755 => x"130101ff",
        1756 => x"b7070020",
        1757 => x"23248100",
        1758 => x"23261100",
        1759 => x"93870709",
        1760 => x"13040500",
        1761 => x"6384f500",
        1762 => x"ef109012",
        1763 => x"83258400",
        1764 => x"9387818f",
        1765 => x"6386f500",
        1766 => x"13050400",
        1767 => x"ef105011",
        1768 => x"8325c400",
        1769 => x"93870196",
        1770 => x"638cf500",
        1771 => x"13050400",
        1772 => x"03248100",
        1773 => x"8320c100",
        1774 => x"13010101",
        1775 => x"6f10500f",
        1776 => x"8320c100",
        1777 => x"03248100",
        1778 => x"13010101",
        1779 => x"67800000",
        1780 => x"b7270000",
        1781 => x"37050020",
        1782 => x"130101ff",
        1783 => x"938707b5",
        1784 => x"13060000",
        1785 => x"93054000",
        1786 => x"13050509",
        1787 => x"23261100",
        1788 => x"23a0f188",
        1789 => x"eff05fed",
        1790 => x"13061000",
        1791 => x"93059000",
        1792 => x"1385818f",
        1793 => x"eff05fec",
        1794 => x"8320c100",
        1795 => x"13062000",
        1796 => x"93052001",
        1797 => x"13850196",
        1798 => x"13010101",
        1799 => x"6ff0dfea",
        1800 => x"13050000",
        1801 => x"67800000",
        1802 => x"83a70188",
        1803 => x"130101ff",
        1804 => x"23202101",
        1805 => x"23261100",
        1806 => x"23248100",
        1807 => x"23229100",
        1808 => x"13090500",
        1809 => x"63940700",
        1810 => x"eff09ff8",
        1811 => x"93848181",
        1812 => x"03a48400",
        1813 => x"83a74400",
        1814 => x"9387f7ff",
        1815 => x"63d80702",
        1816 => x"83a70400",
        1817 => x"6390070c",
        1818 => x"9305c01a",
        1819 => x"13050900",
        1820 => x"ef001009",
        1821 => x"13040500",
        1822 => x"63140508",
        1823 => x"23a00400",
        1824 => x"9307c000",
        1825 => x"2320f900",
        1826 => x"6f004005",
        1827 => x"0317c400",
        1828 => x"63140706",
        1829 => x"b707ffff",
        1830 => x"93871700",
        1831 => x"23220406",
        1832 => x"23200400",
        1833 => x"23220400",
        1834 => x"23240400",
        1835 => x"2326f400",
        1836 => x"23280400",
        1837 => x"232a0400",
        1838 => x"232c0400",
        1839 => x"13068000",
        1840 => x"93050000",
        1841 => x"1305c405",
        1842 => x"eff08fe6",
        1843 => x"232a0402",
        1844 => x"232c0402",
        1845 => x"23240404",
        1846 => x"23260404",
        1847 => x"8320c100",
        1848 => x"13050400",
        1849 => x"03248100",
        1850 => x"83244100",
        1851 => x"03290100",
        1852 => x"13010101",
        1853 => x"67800000",
        1854 => x"13048406",
        1855 => x"6ff0dff5",
        1856 => x"93074000",
        1857 => x"23200500",
        1858 => x"2322f500",
        1859 => x"1305c500",
        1860 => x"2324a400",
        1861 => x"1306001a",
        1862 => x"93050000",
        1863 => x"eff04fe1",
        1864 => x"23a08400",
        1865 => x"83a40400",
        1866 => x"6ff09ff2",
        1867 => x"83270502",
        1868 => x"639e0700",
        1869 => x"b7270000",
        1870 => x"938787b6",
        1871 => x"2320f502",
        1872 => x"83a70188",
        1873 => x"63940700",
        1874 => x"6ff09fe8",
        1875 => x"67800000",
        1876 => x"67800000",
        1877 => x"67800000",
        1878 => x"b7250000",
        1879 => x"13868181",
        1880 => x"938505ac",
        1881 => x"13050000",
        1882 => x"6f008001",
        1883 => x"b7250000",
        1884 => x"13868181",
        1885 => x"938505c2",
        1886 => x"13050000",
        1887 => x"6f004000",
        1888 => x"130101fd",
        1889 => x"23248102",
        1890 => x"23202103",
        1891 => x"232e3101",
        1892 => x"232c4101",
        1893 => x"23286101",
        1894 => x"23267101",
        1895 => x"23261102",
        1896 => x"23229102",
        1897 => x"232a5101",
        1898 => x"93090500",
        1899 => x"138a0500",
        1900 => x"13040600",
        1901 => x"13090000",
        1902 => x"130b1000",
        1903 => x"930bf0ff",
        1904 => x"83248400",
        1905 => x"832a4400",
        1906 => x"938afaff",
        1907 => x"63de0a02",
        1908 => x"03240400",
        1909 => x"e31604fe",
        1910 => x"8320c102",
        1911 => x"03248102",
        1912 => x"83244102",
        1913 => x"8329c101",
        1914 => x"032a8101",
        1915 => x"832a4101",
        1916 => x"032b0101",
        1917 => x"832bc100",
        1918 => x"13050900",
        1919 => x"03290102",
        1920 => x"13010103",
        1921 => x"67800000",
        1922 => x"83d7c400",
        1923 => x"637efb00",
        1924 => x"8397e400",
        1925 => x"638a7701",
        1926 => x"93850400",
        1927 => x"13850900",
        1928 => x"e7000a00",
        1929 => x"3369a900",
        1930 => x"93848406",
        1931 => x"6ff0dff9",
        1932 => x"130101f6",
        1933 => x"232af108",
        1934 => x"b7070080",
        1935 => x"9387f7ff",
        1936 => x"232ef100",
        1937 => x"2328f100",
        1938 => x"b707ffff",
        1939 => x"2326d108",
        1940 => x"2324b100",
        1941 => x"232cb100",
        1942 => x"93878720",
        1943 => x"9306c108",
        1944 => x"93058100",
        1945 => x"232e1106",
        1946 => x"232af100",
        1947 => x"2328e108",
        1948 => x"232c0109",
        1949 => x"232e1109",
        1950 => x"2322d100",
        1951 => x"ef00d037",
        1952 => x"83278100",
        1953 => x"23800700",
        1954 => x"8320c107",
        1955 => x"1301010a",
        1956 => x"67800000",
        1957 => x"130101f6",
        1958 => x"232af108",
        1959 => x"b7070080",
        1960 => x"9387f7ff",
        1961 => x"232ef100",
        1962 => x"2328f100",
        1963 => x"b707ffff",
        1964 => x"93878720",
        1965 => x"232af100",
        1966 => x"2324a100",
        1967 => x"232ca100",
        1968 => x"03a54187",
        1969 => x"2324c108",
        1970 => x"2326d108",
        1971 => x"13860500",
        1972 => x"93068108",
        1973 => x"93058100",
        1974 => x"232e1106",
        1975 => x"2328e108",
        1976 => x"232c0109",
        1977 => x"232e1109",
        1978 => x"2322d100",
        1979 => x"ef00d030",
        1980 => x"83278100",
        1981 => x"23800700",
        1982 => x"8320c107",
        1983 => x"1301010a",
        1984 => x"67800000",
        1985 => x"130101ff",
        1986 => x"23248100",
        1987 => x"13840500",
        1988 => x"8395e500",
        1989 => x"23261100",
        1990 => x"ef008031",
        1991 => x"63400502",
        1992 => x"83274405",
        1993 => x"b387a700",
        1994 => x"232af404",
        1995 => x"8320c100",
        1996 => x"03248100",
        1997 => x"13010101",
        1998 => x"67800000",
        1999 => x"8357c400",
        2000 => x"37f7ffff",
        2001 => x"1307f7ff",
        2002 => x"b3f7e700",
        2003 => x"2316f400",
        2004 => x"6ff0dffd",
        2005 => x"13050000",
        2006 => x"67800000",
        2007 => x"83d7c500",
        2008 => x"130101fe",
        2009 => x"232c8100",
        2010 => x"232a9100",
        2011 => x"23282101",
        2012 => x"23263101",
        2013 => x"232e1100",
        2014 => x"93f70710",
        2015 => x"93040500",
        2016 => x"13840500",
        2017 => x"13090600",
        2018 => x"93890600",
        2019 => x"638a0700",
        2020 => x"8395e500",
        2021 => x"93062000",
        2022 => x"13060000",
        2023 => x"ef004024",
        2024 => x"8357c400",
        2025 => x"37f7ffff",
        2026 => x"1307f7ff",
        2027 => x"b3f7e700",
        2028 => x"8315e400",
        2029 => x"2316f400",
        2030 => x"03248101",
        2031 => x"8320c101",
        2032 => x"93860900",
        2033 => x"13060900",
        2034 => x"8329c100",
        2035 => x"03290101",
        2036 => x"13850400",
        2037 => x"83244101",
        2038 => x"13010102",
        2039 => x"6f00402a",
        2040 => x"130101ff",
        2041 => x"23248100",
        2042 => x"13840500",
        2043 => x"8395e500",
        2044 => x"23261100",
        2045 => x"ef00c01e",
        2046 => x"1307f0ff",
        2047 => x"8357c400",
        2048 => x"6312e502",
        2049 => x"37f7ffff",
        2050 => x"1307f7ff",
        2051 => x"b3f7e700",
        2052 => x"2316f400",
        2053 => x"8320c100",
        2054 => x"03248100",
        2055 => x"13010101",
        2056 => x"67800000",
        2057 => x"37170000",
        2058 => x"b3e7e700",
        2059 => x"2316f400",
        2060 => x"232aa404",
        2061 => x"6ff01ffe",
        2062 => x"8395e500",
        2063 => x"6f004000",
        2064 => x"130101ff",
        2065 => x"23248100",
        2066 => x"23229100",
        2067 => x"13040500",
        2068 => x"13850500",
        2069 => x"23261100",
        2070 => x"23a20188",
        2071 => x"eff0cfcb",
        2072 => x"9307f0ff",
        2073 => x"6318f500",
        2074 => x"83a74188",
        2075 => x"63840700",
        2076 => x"2320f400",
        2077 => x"8320c100",
        2078 => x"03248100",
        2079 => x"83244100",
        2080 => x"13010101",
        2081 => x"67800000",
        2082 => x"83a74187",
        2083 => x"6388a714",
        2084 => x"8327c501",
        2085 => x"130101fe",
        2086 => x"232c8100",
        2087 => x"232e1100",
        2088 => x"232a9100",
        2089 => x"23282101",
        2090 => x"23263101",
        2091 => x"13040500",
        2092 => x"638a0704",
        2093 => x"83a7c700",
        2094 => x"638c0702",
        2095 => x"93040000",
        2096 => x"13090008",
        2097 => x"8327c401",
        2098 => x"83a7c700",
        2099 => x"b3879700",
        2100 => x"83a50700",
        2101 => x"639c050c",
        2102 => x"93844400",
        2103 => x"e39424ff",
        2104 => x"8327c401",
        2105 => x"13050400",
        2106 => x"83a5c700",
        2107 => x"ef008029",
        2108 => x"8327c401",
        2109 => x"83a50700",
        2110 => x"63860500",
        2111 => x"13050400",
        2112 => x"ef004028",
        2113 => x"83254401",
        2114 => x"63860500",
        2115 => x"13050400",
        2116 => x"ef004027",
        2117 => x"8325c401",
        2118 => x"63860500",
        2119 => x"13050400",
        2120 => x"ef004026",
        2121 => x"83250403",
        2122 => x"63860500",
        2123 => x"13050400",
        2124 => x"ef004025",
        2125 => x"83254403",
        2126 => x"63860500",
        2127 => x"13050400",
        2128 => x"ef004024",
        2129 => x"83258403",
        2130 => x"63860500",
        2131 => x"13050400",
        2132 => x"ef004023",
        2133 => x"83258404",
        2134 => x"63860500",
        2135 => x"13050400",
        2136 => x"ef004022",
        2137 => x"83254404",
        2138 => x"63860500",
        2139 => x"13050400",
        2140 => x"ef004021",
        2141 => x"8325c402",
        2142 => x"63860500",
        2143 => x"13050400",
        2144 => x"ef004020",
        2145 => x"83270402",
        2146 => x"638c0702",
        2147 => x"13050400",
        2148 => x"03248101",
        2149 => x"8320c101",
        2150 => x"83244101",
        2151 => x"03290101",
        2152 => x"8329c100",
        2153 => x"13010102",
        2154 => x"67800700",
        2155 => x"83a90500",
        2156 => x"13050400",
        2157 => x"ef00001d",
        2158 => x"93850900",
        2159 => x"6ff09ff1",
        2160 => x"8320c101",
        2161 => x"03248101",
        2162 => x"83244101",
        2163 => x"03290101",
        2164 => x"8329c100",
        2165 => x"13010102",
        2166 => x"67800000",
        2167 => x"67800000",
        2168 => x"130101ff",
        2169 => x"23248100",
        2170 => x"23229100",
        2171 => x"13040500",
        2172 => x"13850500",
        2173 => x"93050600",
        2174 => x"13860600",
        2175 => x"23261100",
        2176 => x"23a20188",
        2177 => x"eff04fb3",
        2178 => x"9307f0ff",
        2179 => x"6318f500",
        2180 => x"83a74188",
        2181 => x"63840700",
        2182 => x"2320f400",
        2183 => x"8320c100",
        2184 => x"03248100",
        2185 => x"83244100",
        2186 => x"13010101",
        2187 => x"67800000",
        2188 => x"130101ff",
        2189 => x"23248100",
        2190 => x"23229100",
        2191 => x"13040500",
        2192 => x"13850500",
        2193 => x"93050600",
        2194 => x"13860600",
        2195 => x"23261100",
        2196 => x"23a20188",
        2197 => x"eff08fa4",
        2198 => x"9307f0ff",
        2199 => x"6318f500",
        2200 => x"83a74188",
        2201 => x"63840700",
        2202 => x"2320f400",
        2203 => x"8320c100",
        2204 => x"03248100",
        2205 => x"83244100",
        2206 => x"13010101",
        2207 => x"67800000",
        2208 => x"130101ff",
        2209 => x"23248100",
        2210 => x"23229100",
        2211 => x"13040500",
        2212 => x"13850500",
        2213 => x"93050600",
        2214 => x"13860600",
        2215 => x"23261100",
        2216 => x"23a20188",
        2217 => x"eff08f9a",
        2218 => x"9307f0ff",
        2219 => x"6318f500",
        2220 => x"83a74188",
        2221 => x"63840700",
        2222 => x"2320f400",
        2223 => x"8320c100",
        2224 => x"03248100",
        2225 => x"83244100",
        2226 => x"13010101",
        2227 => x"67800000",
        2228 => x"03a54187",
        2229 => x"67800000",
        2230 => x"130101ff",
        2231 => x"23248100",
        2232 => x"23229100",
        2233 => x"37440000",
        2234 => x"b7440000",
        2235 => x"938784b6",
        2236 => x"130484b6",
        2237 => x"3304f440",
        2238 => x"23202101",
        2239 => x"23261100",
        2240 => x"13542440",
        2241 => x"938484b6",
        2242 => x"13090000",
        2243 => x"63108904",
        2244 => x"b7440000",
        2245 => x"37440000",
        2246 => x"938784b6",
        2247 => x"130484b6",
        2248 => x"3304f440",
        2249 => x"13542440",
        2250 => x"938484b6",
        2251 => x"13090000",
        2252 => x"63188902",
        2253 => x"8320c100",
        2254 => x"03248100",
        2255 => x"83244100",
        2256 => x"03290100",
        2257 => x"13010101",
        2258 => x"67800000",
        2259 => x"83a70400",
        2260 => x"13091900",
        2261 => x"93844400",
        2262 => x"e7800700",
        2263 => x"6ff01ffb",
        2264 => x"83a70400",
        2265 => x"13091900",
        2266 => x"93844400",
        2267 => x"e7800700",
        2268 => x"6ff01ffc",
        2269 => x"13860500",
        2270 => x"93050500",
        2271 => x"03a54187",
        2272 => x"6f10401e",
        2273 => x"638a050e",
        2274 => x"83a7c5ff",
        2275 => x"130101fe",
        2276 => x"232c8100",
        2277 => x"232e1100",
        2278 => x"1384c5ff",
        2279 => x"63d40700",
        2280 => x"3304f400",
        2281 => x"2326a100",
        2282 => x"ef008031",
        2283 => x"83a7c188",
        2284 => x"0325c100",
        2285 => x"639e0700",
        2286 => x"23220400",
        2287 => x"23a68188",
        2288 => x"03248101",
        2289 => x"8320c101",
        2290 => x"13010102",
        2291 => x"6f00802f",
        2292 => x"6374f402",
        2293 => x"03260400",
        2294 => x"b306c400",
        2295 => x"639ad700",
        2296 => x"83a60700",
        2297 => x"83a74700",
        2298 => x"b386c600",
        2299 => x"2320d400",
        2300 => x"2322f400",
        2301 => x"6ff09ffc",
        2302 => x"13870700",
        2303 => x"83a74700",
        2304 => x"63840700",
        2305 => x"e37af4fe",
        2306 => x"83260700",
        2307 => x"3306d700",
        2308 => x"63188602",
        2309 => x"03260400",
        2310 => x"b386c600",
        2311 => x"2320d700",
        2312 => x"3306d700",
        2313 => x"e39ec7f8",
        2314 => x"03a60700",
        2315 => x"83a74700",
        2316 => x"b306d600",
        2317 => x"2320d700",
        2318 => x"2322f700",
        2319 => x"6ff05ff8",
        2320 => x"6378c400",
        2321 => x"9307c000",
        2322 => x"2320f500",
        2323 => x"6ff05ff7",
        2324 => x"03260400",
        2325 => x"b306c400",
        2326 => x"639ad700",
        2327 => x"83a60700",
        2328 => x"83a74700",
        2329 => x"b386c600",
        2330 => x"2320d400",
        2331 => x"2322f400",
        2332 => x"23228700",
        2333 => x"6ff0dff4",
        2334 => x"67800000",
        2335 => x"130101ff",
        2336 => x"23202101",
        2337 => x"83a78188",
        2338 => x"23248100",
        2339 => x"23229100",
        2340 => x"23261100",
        2341 => x"93040500",
        2342 => x"13840500",
        2343 => x"63980700",
        2344 => x"93050000",
        2345 => x"ef10c010",
        2346 => x"23a4a188",
        2347 => x"93050400",
        2348 => x"13850400",
        2349 => x"ef10c00f",
        2350 => x"1309f0ff",
        2351 => x"63122503",
        2352 => x"1304f0ff",
        2353 => x"8320c100",
        2354 => x"13050400",
        2355 => x"03248100",
        2356 => x"83244100",
        2357 => x"03290100",
        2358 => x"13010101",
        2359 => x"67800000",
        2360 => x"13043500",
        2361 => x"1374c4ff",
        2362 => x"e30e85fc",
        2363 => x"b305a440",
        2364 => x"13850400",
        2365 => x"ef10c00b",
        2366 => x"e31625fd",
        2367 => x"6ff05ffc",
        2368 => x"130101fe",
        2369 => x"232a9100",
        2370 => x"93843500",
        2371 => x"93f4c4ff",
        2372 => x"23282101",
        2373 => x"232e1100",
        2374 => x"232c8100",
        2375 => x"23263101",
        2376 => x"23244101",
        2377 => x"93848400",
        2378 => x"9307c000",
        2379 => x"13090500",
        2380 => x"63f0f40a",
        2381 => x"9304c000",
        2382 => x"63eeb408",
        2383 => x"13050900",
        2384 => x"ef000018",
        2385 => x"83a7c188",
        2386 => x"13840700",
        2387 => x"631a040a",
        2388 => x"93850400",
        2389 => x"13050900",
        2390 => x"eff05ff2",
        2391 => x"9307f0ff",
        2392 => x"13040500",
        2393 => x"6316f514",
        2394 => x"03a4c188",
        2395 => x"93070400",
        2396 => x"639c0710",
        2397 => x"63040412",
        2398 => x"032a0400",
        2399 => x"93050000",
        2400 => x"13050900",
        2401 => x"330a4401",
        2402 => x"ef108002",
        2403 => x"6318aa10",
        2404 => x"83270400",
        2405 => x"13050900",
        2406 => x"b384f440",
        2407 => x"93850400",
        2408 => x"eff0dfed",
        2409 => x"9307f0ff",
        2410 => x"630af50e",
        2411 => x"83270400",
        2412 => x"b3879700",
        2413 => x"2320f400",
        2414 => x"83a7c188",
        2415 => x"638e070e",
        2416 => x"03a74700",
        2417 => x"6318870c",
        2418 => x"23a20700",
        2419 => x"6f004006",
        2420 => x"e3d404f6",
        2421 => x"9307c000",
        2422 => x"2320f900",
        2423 => x"13050000",
        2424 => x"8320c101",
        2425 => x"03248101",
        2426 => x"83244101",
        2427 => x"03290101",
        2428 => x"8329c100",
        2429 => x"032a8100",
        2430 => x"13010102",
        2431 => x"67800000",
        2432 => x"83260400",
        2433 => x"b3869640",
        2434 => x"63ca0606",
        2435 => x"1307b000",
        2436 => x"637ad704",
        2437 => x"23209400",
        2438 => x"33079400",
        2439 => x"63908704",
        2440 => x"23a6e188",
        2441 => x"83274400",
        2442 => x"2320d700",
        2443 => x"2322f700",
        2444 => x"13050900",
        2445 => x"ef000009",
        2446 => x"1305b400",
        2447 => x"93074400",
        2448 => x"137585ff",
        2449 => x"3307f540",
        2450 => x"e30cf5f8",
        2451 => x"3304e400",
        2452 => x"b387a740",
        2453 => x"2320f400",
        2454 => x"6ff09ff8",
        2455 => x"23a2e700",
        2456 => x"6ff05ffc",
        2457 => x"03274400",
        2458 => x"63968700",
        2459 => x"23a6e188",
        2460 => x"6ff01ffc",
        2461 => x"23a2e700",
        2462 => x"6ff09ffb",
        2463 => x"93070400",
        2464 => x"03244400",
        2465 => x"6ff09fec",
        2466 => x"13840700",
        2467 => x"83a74700",
        2468 => x"6ff01fee",
        2469 => x"93070700",
        2470 => x"6ff05ff2",
        2471 => x"9307c000",
        2472 => x"2320f900",
        2473 => x"13050900",
        2474 => x"ef00c001",
        2475 => x"6ff01ff3",
        2476 => x"23209500",
        2477 => x"6ff0dff7",
        2478 => x"23220000",
        2479 => x"73001000",
        2480 => x"67800000",
        2481 => x"67800000",
        2482 => x"130101fe",
        2483 => x"23282101",
        2484 => x"03a98500",
        2485 => x"232c8100",
        2486 => x"23263101",
        2487 => x"23225101",
        2488 => x"23206101",
        2489 => x"232e1100",
        2490 => x"232a9100",
        2491 => x"23244101",
        2492 => x"83aa0500",
        2493 => x"13840500",
        2494 => x"130b0600",
        2495 => x"93890600",
        2496 => x"63ec2609",
        2497 => x"8397c500",
        2498 => x"13f70748",
        2499 => x"63040708",
        2500 => x"03274401",
        2501 => x"93043000",
        2502 => x"83a50501",
        2503 => x"b384e402",
        2504 => x"13072000",
        2505 => x"b38aba40",
        2506 => x"130a0500",
        2507 => x"b3c4e402",
        2508 => x"13871600",
        2509 => x"33075701",
        2510 => x"63f4e400",
        2511 => x"93040700",
        2512 => x"93f70740",
        2513 => x"6386070a",
        2514 => x"93850400",
        2515 => x"13050a00",
        2516 => x"eff01fdb",
        2517 => x"13090500",
        2518 => x"630c050a",
        2519 => x"83250401",
        2520 => x"13860a00",
        2521 => x"efe09fbe",
        2522 => x"8357c400",
        2523 => x"93f7f7b7",
        2524 => x"93e70708",
        2525 => x"2316f400",
        2526 => x"23282401",
        2527 => x"232a9400",
        2528 => x"33095901",
        2529 => x"b3845441",
        2530 => x"23202401",
        2531 => x"23249400",
        2532 => x"13890900",
        2533 => x"63f42901",
        2534 => x"13890900",
        2535 => x"03250400",
        2536 => x"13060900",
        2537 => x"93050b00",
        2538 => x"efe09fbc",
        2539 => x"83278400",
        2540 => x"13050000",
        2541 => x"b3872741",
        2542 => x"2324f400",
        2543 => x"83270400",
        2544 => x"b3872701",
        2545 => x"2320f400",
        2546 => x"8320c101",
        2547 => x"03248101",
        2548 => x"83244101",
        2549 => x"03290101",
        2550 => x"8329c100",
        2551 => x"032a8100",
        2552 => x"832a4100",
        2553 => x"032b0100",
        2554 => x"13010102",
        2555 => x"67800000",
        2556 => x"13860400",
        2557 => x"13050a00",
        2558 => x"ef001060",
        2559 => x"13090500",
        2560 => x"e31c05f6",
        2561 => x"83250401",
        2562 => x"13050a00",
        2563 => x"eff09fb7",
        2564 => x"9307c000",
        2565 => x"2320fa00",
        2566 => x"8357c400",
        2567 => x"1305f0ff",
        2568 => x"93e70704",
        2569 => x"2316f400",
        2570 => x"6ff01ffa",
        2571 => x"83278600",
        2572 => x"130101fd",
        2573 => x"232e3101",
        2574 => x"23267101",
        2575 => x"23261102",
        2576 => x"23248102",
        2577 => x"23229102",
        2578 => x"23202103",
        2579 => x"232c4101",
        2580 => x"232a5101",
        2581 => x"23286101",
        2582 => x"23248101",
        2583 => x"23229101",
        2584 => x"2320a101",
        2585 => x"832b0600",
        2586 => x"93090600",
        2587 => x"63980712",
        2588 => x"13050000",
        2589 => x"8320c102",
        2590 => x"03248102",
        2591 => x"23a20900",
        2592 => x"83244102",
        2593 => x"03290102",
        2594 => x"8329c101",
        2595 => x"032a8101",
        2596 => x"832a4101",
        2597 => x"032b0101",
        2598 => x"832bc100",
        2599 => x"032c8100",
        2600 => x"832c4100",
        2601 => x"032d0100",
        2602 => x"13010103",
        2603 => x"67800000",
        2604 => x"03ab0b00",
        2605 => x"03ad4b00",
        2606 => x"938b8b00",
        2607 => x"03298400",
        2608 => x"832a0400",
        2609 => x"e3060dfe",
        2610 => x"63642d09",
        2611 => x"8317c400",
        2612 => x"13f70748",
        2613 => x"63020708",
        2614 => x"83244401",
        2615 => x"83250401",
        2616 => x"b3049c02",
        2617 => x"b38aba40",
        2618 => x"13871a00",
        2619 => x"3307a701",
        2620 => x"b3c49403",
        2621 => x"63f4e400",
        2622 => x"93040700",
        2623 => x"93f70740",
        2624 => x"638c070a",
        2625 => x"93850400",
        2626 => x"13050a00",
        2627 => x"eff05fbf",
        2628 => x"13090500",
        2629 => x"6302050c",
        2630 => x"83250401",
        2631 => x"13860a00",
        2632 => x"efe0dfa2",
        2633 => x"8357c400",
        2634 => x"93f7f7b7",
        2635 => x"93e70708",
        2636 => x"2316f400",
        2637 => x"23282401",
        2638 => x"232a9400",
        2639 => x"33095901",
        2640 => x"b3845441",
        2641 => x"23202401",
        2642 => x"23249400",
        2643 => x"13090d00",
        2644 => x"63742d01",
        2645 => x"13090d00",
        2646 => x"03250400",
        2647 => x"93050b00",
        2648 => x"13060900",
        2649 => x"efe0dfa0",
        2650 => x"83278400",
        2651 => x"330bab01",
        2652 => x"b3872741",
        2653 => x"2324f400",
        2654 => x"83270400",
        2655 => x"b3872701",
        2656 => x"2320f400",
        2657 => x"83a78900",
        2658 => x"b387a741",
        2659 => x"23a4f900",
        2660 => x"e38007ee",
        2661 => x"130d0000",
        2662 => x"6ff05ff2",
        2663 => x"130a0500",
        2664 => x"13840500",
        2665 => x"130b0000",
        2666 => x"130d0000",
        2667 => x"130c3000",
        2668 => x"930c2000",
        2669 => x"6ff09ff0",
        2670 => x"13860400",
        2671 => x"13050a00",
        2672 => x"ef009043",
        2673 => x"13090500",
        2674 => x"e31605f6",
        2675 => x"83250401",
        2676 => x"13050a00",
        2677 => x"eff01f9b",
        2678 => x"9307c000",
        2679 => x"2320fa00",
        2680 => x"8357c400",
        2681 => x"1305f0ff",
        2682 => x"93e70704",
        2683 => x"2316f400",
        2684 => x"23a40900",
        2685 => x"6ff01fe8",
        2686 => x"83d7c500",
        2687 => x"130101f5",
        2688 => x"2324810a",
        2689 => x"2322910a",
        2690 => x"2320210b",
        2691 => x"232c4109",
        2692 => x"2326110a",
        2693 => x"232e3109",
        2694 => x"232a5109",
        2695 => x"23286109",
        2696 => x"23267109",
        2697 => x"23248109",
        2698 => x"23229109",
        2699 => x"2320a109",
        2700 => x"232eb107",
        2701 => x"93f70708",
        2702 => x"130a0500",
        2703 => x"13890500",
        2704 => x"93040600",
        2705 => x"13840600",
        2706 => x"63880706",
        2707 => x"83a70501",
        2708 => x"63940706",
        2709 => x"93050004",
        2710 => x"eff09faa",
        2711 => x"2320a900",
        2712 => x"2328a900",
        2713 => x"63160504",
        2714 => x"9307c000",
        2715 => x"2320fa00",
        2716 => x"1305f0ff",
        2717 => x"8320c10a",
        2718 => x"0324810a",
        2719 => x"8324410a",
        2720 => x"0329010a",
        2721 => x"8329c109",
        2722 => x"032a8109",
        2723 => x"832a4109",
        2724 => x"032b0109",
        2725 => x"832bc108",
        2726 => x"032c8108",
        2727 => x"832c4108",
        2728 => x"032d0108",
        2729 => x"832dc107",
        2730 => x"1301010b",
        2731 => x"67800000",
        2732 => x"93070004",
        2733 => x"232af900",
        2734 => x"93070002",
        2735 => x"a304f102",
        2736 => x"93070003",
        2737 => x"23220102",
        2738 => x"2305f102",
        2739 => x"23268100",
        2740 => x"930c5002",
        2741 => x"374b0000",
        2742 => x"b74b0000",
        2743 => x"374d0000",
        2744 => x"372c0000",
        2745 => x"930a0000",
        2746 => x"13840400",
        2747 => x"83470400",
        2748 => x"63840700",
        2749 => x"639c970d",
        2750 => x"b30d9440",
        2751 => x"63069402",
        2752 => x"93860d00",
        2753 => x"13860400",
        2754 => x"93050900",
        2755 => x"13050a00",
        2756 => x"eff09fbb",
        2757 => x"9307f0ff",
        2758 => x"6304f524",
        2759 => x"83274102",
        2760 => x"b387b701",
        2761 => x"2322f102",
        2762 => x"83470400",
        2763 => x"638a0722",
        2764 => x"9307f0ff",
        2765 => x"93041400",
        2766 => x"23280100",
        2767 => x"232e0100",
        2768 => x"232af100",
        2769 => x"232c0100",
        2770 => x"a3090104",
        2771 => x"23240106",
        2772 => x"930d1000",
        2773 => x"83c50400",
        2774 => x"13065000",
        2775 => x"13054bad",
        2776 => x"ef00101e",
        2777 => x"83270101",
        2778 => x"13841400",
        2779 => x"63140506",
        2780 => x"13f70701",
        2781 => x"63060700",
        2782 => x"13070002",
        2783 => x"a309e104",
        2784 => x"13f78700",
        2785 => x"63060700",
        2786 => x"1307b002",
        2787 => x"a309e104",
        2788 => x"83c60400",
        2789 => x"1307a002",
        2790 => x"638ce604",
        2791 => x"8327c101",
        2792 => x"13840400",
        2793 => x"93060000",
        2794 => x"13069000",
        2795 => x"1305a000",
        2796 => x"03470400",
        2797 => x"93051400",
        2798 => x"130707fd",
        2799 => x"637ee608",
        2800 => x"63840604",
        2801 => x"232ef100",
        2802 => x"6f000004",
        2803 => x"13041400",
        2804 => x"6ff0dff1",
        2805 => x"13074bad",
        2806 => x"3305e540",
        2807 => x"3395ad00",
        2808 => x"b3e7a700",
        2809 => x"2328f100",
        2810 => x"93040400",
        2811 => x"6ff09ff6",
        2812 => x"0327c100",
        2813 => x"93064700",
        2814 => x"03270700",
        2815 => x"2326d100",
        2816 => x"63420704",
        2817 => x"232ee100",
        2818 => x"03470400",
        2819 => x"9307e002",
        2820 => x"6314f708",
        2821 => x"03471400",
        2822 => x"9307a002",
        2823 => x"6318f704",
        2824 => x"8327c100",
        2825 => x"13042400",
        2826 => x"13874700",
        2827 => x"83a70700",
        2828 => x"2326e100",
        2829 => x"63d40700",
        2830 => x"9307f0ff",
        2831 => x"232af100",
        2832 => x"6f008005",
        2833 => x"3307e040",
        2834 => x"93e72700",
        2835 => x"232ee100",
        2836 => x"2328f100",
        2837 => x"6ff05ffb",
        2838 => x"b387a702",
        2839 => x"13840500",
        2840 => x"93061000",
        2841 => x"b387e700",
        2842 => x"6ff09ff4",
        2843 => x"13041400",
        2844 => x"232a0100",
        2845 => x"93060000",
        2846 => x"93070000",
        2847 => x"13069000",
        2848 => x"1305a000",
        2849 => x"03470400",
        2850 => x"93051400",
        2851 => x"130707fd",
        2852 => x"6372e608",
        2853 => x"e39406fa",
        2854 => x"83450400",
        2855 => x"13063000",
        2856 => x"1385cbad",
        2857 => x"ef00d009",
        2858 => x"63020502",
        2859 => x"9387cbad",
        2860 => x"3305f540",
        2861 => x"83270101",
        2862 => x"13070004",
        2863 => x"3317a700",
        2864 => x"b3e7e700",
        2865 => x"13041400",
        2866 => x"2328f100",
        2867 => x"83450400",
        2868 => x"13066000",
        2869 => x"13050dae",
        2870 => x"93041400",
        2871 => x"2304b102",
        2872 => x"ef001006",
        2873 => x"63080508",
        2874 => x"63980a04",
        2875 => x"03270101",
        2876 => x"8327c100",
        2877 => x"13770710",
        2878 => x"63080702",
        2879 => x"93874700",
        2880 => x"2326f100",
        2881 => x"83274102",
        2882 => x"b3873701",
        2883 => x"2322f102",
        2884 => x"6ff09fdd",
        2885 => x"b387a702",
        2886 => x"13840500",
        2887 => x"93061000",
        2888 => x"b387e700",
        2889 => x"6ff01ff6",
        2890 => x"93877700",
        2891 => x"93f787ff",
        2892 => x"93878700",
        2893 => x"6ff0dffc",
        2894 => x"1307c100",
        2895 => x"93068c6c",
        2896 => x"13060900",
        2897 => x"93050101",
        2898 => x"13050a00",
        2899 => x"97000000",
        2900 => x"e7000000",
        2901 => x"9307f0ff",
        2902 => x"93090500",
        2903 => x"e314f5fa",
        2904 => x"8357c900",
        2905 => x"93f70704",
        2906 => x"e39407d0",
        2907 => x"03254102",
        2908 => x"6ff05fd0",
        2909 => x"1307c100",
        2910 => x"93068c6c",
        2911 => x"13060900",
        2912 => x"93050101",
        2913 => x"13050a00",
        2914 => x"ef00801b",
        2915 => x"6ff09ffc",
        2916 => x"130101fd",
        2917 => x"232a5101",
        2918 => x"83a70501",
        2919 => x"930a0700",
        2920 => x"03a78500",
        2921 => x"23248102",
        2922 => x"23202103",
        2923 => x"232e3101",
        2924 => x"232c4101",
        2925 => x"23261102",
        2926 => x"23229102",
        2927 => x"23286101",
        2928 => x"23267101",
        2929 => x"93090500",
        2930 => x"13840500",
        2931 => x"13090600",
        2932 => x"138a0600",
        2933 => x"63d4e700",
        2934 => x"93070700",
        2935 => x"2320f900",
        2936 => x"03473404",
        2937 => x"63060700",
        2938 => x"93871700",
        2939 => x"2320f900",
        2940 => x"83270400",
        2941 => x"93f70702",
        2942 => x"63880700",
        2943 => x"83270900",
        2944 => x"93872700",
        2945 => x"2320f900",
        2946 => x"83240400",
        2947 => x"93f46400",
        2948 => x"639e0400",
        2949 => x"130b9401",
        2950 => x"930bf0ff",
        2951 => x"8327c400",
        2952 => x"03270900",
        2953 => x"b387e740",
        2954 => x"63c2f408",
        2955 => x"83473404",
        2956 => x"b336f000",
        2957 => x"83270400",
        2958 => x"93f70702",
        2959 => x"6390070c",
        2960 => x"13063404",
        2961 => x"93050a00",
        2962 => x"13850900",
        2963 => x"e7800a00",
        2964 => x"9307f0ff",
        2965 => x"6308f506",
        2966 => x"83270400",
        2967 => x"13074000",
        2968 => x"93040000",
        2969 => x"93f76700",
        2970 => x"639ce700",
        2971 => x"8324c400",
        2972 => x"83270900",
        2973 => x"b384f440",
        2974 => x"63d40400",
        2975 => x"93040000",
        2976 => x"83278400",
        2977 => x"03270401",
        2978 => x"6356f700",
        2979 => x"b387e740",
        2980 => x"b384f400",
        2981 => x"13090000",
        2982 => x"1304a401",
        2983 => x"130bf0ff",
        2984 => x"63902409",
        2985 => x"13050000",
        2986 => x"6f000002",
        2987 => x"93061000",
        2988 => x"13060b00",
        2989 => x"93050a00",
        2990 => x"13850900",
        2991 => x"e7800a00",
        2992 => x"631a7503",
        2993 => x"1305f0ff",
        2994 => x"8320c102",
        2995 => x"03248102",
        2996 => x"83244102",
        2997 => x"03290102",
        2998 => x"8329c101",
        2999 => x"032a8101",
        3000 => x"832a4101",
        3001 => x"032b0101",
        3002 => x"832bc100",
        3003 => x"13010103",
        3004 => x"67800000",
        3005 => x"93841400",
        3006 => x"6ff05ff2",
        3007 => x"3307d400",
        3008 => x"13060003",
        3009 => x"a301c704",
        3010 => x"03475404",
        3011 => x"93871600",
        3012 => x"b307f400",
        3013 => x"93862600",
        3014 => x"a381e704",
        3015 => x"6ff05ff2",
        3016 => x"93061000",
        3017 => x"13060400",
        3018 => x"93050a00",
        3019 => x"13850900",
        3020 => x"e7800a00",
        3021 => x"e30865f9",
        3022 => x"13091900",
        3023 => x"6ff05ff6",
        3024 => x"130101fd",
        3025 => x"23248102",
        3026 => x"23202103",
        3027 => x"232e3101",
        3028 => x"232c4101",
        3029 => x"23261102",
        3030 => x"23229102",
        3031 => x"232a5101",
        3032 => x"23286101",
        3033 => x"138a0600",
        3034 => x"83c68501",
        3035 => x"93078007",
        3036 => x"13090500",
        3037 => x"13840500",
        3038 => x"93090600",
        3039 => x"63eed700",
        3040 => x"93072006",
        3041 => x"13863504",
        3042 => x"63eed700",
        3043 => x"63840628",
        3044 => x"93078005",
        3045 => x"6380f622",
        3046 => x"93042404",
        3047 => x"2301d404",
        3048 => x"6f004004",
        3049 => x"9387d6f9",
        3050 => x"93f7f70f",
        3051 => x"93055001",
        3052 => x"e3e4f5fe",
        3053 => x"b7450000",
        3054 => x"93972700",
        3055 => x"938505b1",
        3056 => x"b387b700",
        3057 => x"83a70700",
        3058 => x"67800700",
        3059 => x"83270700",
        3060 => x"93042404",
        3061 => x"93864700",
        3062 => x"83a70700",
        3063 => x"2320d700",
        3064 => x"2301f404",
        3065 => x"93071000",
        3066 => x"6f008026",
        3067 => x"83270400",
        3068 => x"03250700",
        3069 => x"93f60708",
        3070 => x"93054500",
        3071 => x"63860602",
        3072 => x"83270500",
        3073 => x"2320b700",
        3074 => x"37480000",
        3075 => x"63d80700",
        3076 => x"1307d002",
        3077 => x"b307f040",
        3078 => x"a301e404",
        3079 => x"130888ae",
        3080 => x"1307a000",
        3081 => x"6f004006",
        3082 => x"93f60704",
        3083 => x"83270500",
        3084 => x"2320b700",
        3085 => x"e38a06fc",
        3086 => x"93970701",
        3087 => x"93d70741",
        3088 => x"6ff09ffc",
        3089 => x"03250400",
        3090 => x"83250700",
        3091 => x"13780508",
        3092 => x"83a70500",
        3093 => x"93854500",
        3094 => x"631a0800",
        3095 => x"13750504",
        3096 => x"63060500",
        3097 => x"93970701",
        3098 => x"93d70701",
        3099 => x"2320b700",
        3100 => x"37480000",
        3101 => x"1307f006",
        3102 => x"130888ae",
        3103 => x"639ae614",
        3104 => x"13078000",
        3105 => x"a3010404",
        3106 => x"83264400",
        3107 => x"2324d400",
        3108 => x"63ce0600",
        3109 => x"83250400",
        3110 => x"b3e6d700",
        3111 => x"93040600",
        3112 => x"93f5b5ff",
        3113 => x"2320b400",
        3114 => x"63840602",
        3115 => x"93040600",
        3116 => x"b3f6e702",
        3117 => x"9384f4ff",
        3118 => x"b306d800",
        3119 => x"83c60600",
        3120 => x"2380d400",
        3121 => x"93860700",
        3122 => x"b3d7e702",
        3123 => x"e3f2e6fe",
        3124 => x"93078000",
        3125 => x"6314f702",
        3126 => x"83270400",
        3127 => x"93f71700",
        3128 => x"638e0700",
        3129 => x"03274400",
        3130 => x"83270401",
        3131 => x"63c8e700",
        3132 => x"93070003",
        3133 => x"a38ff4fe",
        3134 => x"9384f4ff",
        3135 => x"33069640",
        3136 => x"2328c400",
        3137 => x"13070a00",
        3138 => x"93860900",
        3139 => x"1306c100",
        3140 => x"93050400",
        3141 => x"13050900",
        3142 => x"eff09fc7",
        3143 => x"930af0ff",
        3144 => x"631e5513",
        3145 => x"1305f0ff",
        3146 => x"8320c102",
        3147 => x"03248102",
        3148 => x"83244102",
        3149 => x"03290102",
        3150 => x"8329c101",
        3151 => x"032a8101",
        3152 => x"832a4101",
        3153 => x"032b0101",
        3154 => x"13010103",
        3155 => x"67800000",
        3156 => x"83270400",
        3157 => x"93e70702",
        3158 => x"2320f400",
        3159 => x"37480000",
        3160 => x"93068007",
        3161 => x"1308c8af",
        3162 => x"a302d404",
        3163 => x"83260400",
        3164 => x"83250700",
        3165 => x"13f50608",
        3166 => x"83a70500",
        3167 => x"93854500",
        3168 => x"631a0500",
        3169 => x"13f50604",
        3170 => x"63060500",
        3171 => x"93970701",
        3172 => x"93d70701",
        3173 => x"2320b700",
        3174 => x"13f71600",
        3175 => x"63060700",
        3176 => x"93e60602",
        3177 => x"2320d400",
        3178 => x"638c0700",
        3179 => x"13070001",
        3180 => x"6ff05fed",
        3181 => x"37480000",
        3182 => x"130888ae",
        3183 => x"6ff0dffa",
        3184 => x"03270400",
        3185 => x"1377f7fd",
        3186 => x"2320e400",
        3187 => x"6ff01ffe",
        3188 => x"1307a000",
        3189 => x"6ff01feb",
        3190 => x"83260400",
        3191 => x"83270700",
        3192 => x"83254401",
        3193 => x"13f80608",
        3194 => x"13854700",
        3195 => x"630a0800",
        3196 => x"2320a700",
        3197 => x"83a70700",
        3198 => x"23a0b700",
        3199 => x"6f008001",
        3200 => x"2320a700",
        3201 => x"93f60604",
        3202 => x"83a70700",
        3203 => x"e38606fe",
        3204 => x"2390b700",
        3205 => x"23280400",
        3206 => x"93040600",
        3207 => x"6ff09fee",
        3208 => x"83270700",
        3209 => x"03264400",
        3210 => x"93050000",
        3211 => x"93864700",
        3212 => x"2320d700",
        3213 => x"83a40700",
        3214 => x"13850400",
        3215 => x"ef004030",
        3216 => x"63060500",
        3217 => x"33059540",
        3218 => x"2322a400",
        3219 => x"83274400",
        3220 => x"2328f400",
        3221 => x"a3010404",
        3222 => x"6ff0dfea",
        3223 => x"83260401",
        3224 => x"13860400",
        3225 => x"93850900",
        3226 => x"13050900",
        3227 => x"e7000a00",
        3228 => x"e30a55eb",
        3229 => x"83270400",
        3230 => x"93f72700",
        3231 => x"63940704",
        3232 => x"8327c100",
        3233 => x"0325c400",
        3234 => x"e350f5ea",
        3235 => x"13850700",
        3236 => x"6ff09fe9",
        3237 => x"93061000",
        3238 => x"13860a00",
        3239 => x"93850900",
        3240 => x"13050900",
        3241 => x"e7000a00",
        3242 => x"e30e65e7",
        3243 => x"93841400",
        3244 => x"8327c400",
        3245 => x"0327c100",
        3246 => x"b387e740",
        3247 => x"e3ccf4fc",
        3248 => x"6ff01ffc",
        3249 => x"93040000",
        3250 => x"930a9401",
        3251 => x"130bf0ff",
        3252 => x"6ff01ffe",
        3253 => x"8397c500",
        3254 => x"130101fe",
        3255 => x"232c8100",
        3256 => x"232a9100",
        3257 => x"232e1100",
        3258 => x"23282101",
        3259 => x"23263101",
        3260 => x"13f78700",
        3261 => x"93040500",
        3262 => x"13840500",
        3263 => x"631a0712",
        3264 => x"03a74500",
        3265 => x"6346e000",
        3266 => x"03a70504",
        3267 => x"6356e010",
        3268 => x"0327c402",
        3269 => x"63020710",
        3270 => x"03a90400",
        3271 => x"93963701",
        3272 => x"23a00400",
        3273 => x"83250402",
        3274 => x"63dc060a",
        3275 => x"03264405",
        3276 => x"8357c400",
        3277 => x"93f74700",
        3278 => x"638e0700",
        3279 => x"83274400",
        3280 => x"3306f640",
        3281 => x"83274403",
        3282 => x"63860700",
        3283 => x"83270404",
        3284 => x"3306f640",
        3285 => x"8327c402",
        3286 => x"83250402",
        3287 => x"93060000",
        3288 => x"13850400",
        3289 => x"e7800700",
        3290 => x"1307f0ff",
        3291 => x"8357c400",
        3292 => x"6312e502",
        3293 => x"83a60400",
        3294 => x"1307d001",
        3295 => x"6362d70a",
        3296 => x"37074020",
        3297 => x"13071700",
        3298 => x"3357d700",
        3299 => x"13771700",
        3300 => x"63080708",
        3301 => x"03270401",
        3302 => x"23220400",
        3303 => x"2320e400",
        3304 => x"13973701",
        3305 => x"635c0700",
        3306 => x"9307f0ff",
        3307 => x"6316f500",
        3308 => x"83a70400",
        3309 => x"63940700",
        3310 => x"232aa404",
        3311 => x"83254403",
        3312 => x"23a02401",
        3313 => x"638a0504",
        3314 => x"93074404",
        3315 => x"6386f500",
        3316 => x"13850400",
        3317 => x"efe01ffb",
        3318 => x"232a0402",
        3319 => x"6f00c003",
        3320 => x"13060000",
        3321 => x"93061000",
        3322 => x"13850400",
        3323 => x"e7000700",
        3324 => x"9307f0ff",
        3325 => x"13060500",
        3326 => x"e31cf5f2",
        3327 => x"83a70400",
        3328 => x"e38807f2",
        3329 => x"1307d001",
        3330 => x"6386e700",
        3331 => x"13076001",
        3332 => x"6394e706",
        3333 => x"23a02401",
        3334 => x"13050000",
        3335 => x"6f00c006",
        3336 => x"93e70704",
        3337 => x"93970701",
        3338 => x"93d70741",
        3339 => x"6f004005",
        3340 => x"83a90501",
        3341 => x"e38209fe",
        3342 => x"03a90500",
        3343 => x"93f73700",
        3344 => x"23a03501",
        3345 => x"33093941",
        3346 => x"13070000",
        3347 => x"63940700",
        3348 => x"03a74501",
        3349 => x"2324e400",
        3350 => x"e35020fd",
        3351 => x"83278402",
        3352 => x"83250402",
        3353 => x"93060900",
        3354 => x"13860900",
        3355 => x"13850400",
        3356 => x"e7800700",
        3357 => x"6348a002",
        3358 => x"8317c400",
        3359 => x"93e70704",
        3360 => x"2316f400",
        3361 => x"1305f0ff",
        3362 => x"8320c101",
        3363 => x"03248101",
        3364 => x"83244101",
        3365 => x"03290101",
        3366 => x"8329c100",
        3367 => x"13010102",
        3368 => x"67800000",
        3369 => x"b389a900",
        3370 => x"3309a940",
        3371 => x"6ff0dffa",
        3372 => x"83a70501",
        3373 => x"638e0704",
        3374 => x"130101fe",
        3375 => x"232c8100",
        3376 => x"232e1100",
        3377 => x"13040500",
        3378 => x"630c0500",
        3379 => x"83270502",
        3380 => x"63980700",
        3381 => x"2326b100",
        3382 => x"efe05f85",
        3383 => x"8325c100",
        3384 => x"8397c500",
        3385 => x"638c0700",
        3386 => x"13050400",
        3387 => x"03248101",
        3388 => x"8320c101",
        3389 => x"13010102",
        3390 => x"6ff0dfdd",
        3391 => x"8320c101",
        3392 => x"03248101",
        3393 => x"13050000",
        3394 => x"13010102",
        3395 => x"67800000",
        3396 => x"13050000",
        3397 => x"67800000",
        3398 => x"93050500",
        3399 => x"631e0500",
        3400 => x"b7350000",
        3401 => x"37050020",
        3402 => x"13868181",
        3403 => x"9385054b",
        3404 => x"13054502",
        3405 => x"6fe0df84",
        3406 => x"03a54187",
        3407 => x"6ff05ff7",
        3408 => x"93f5f50f",
        3409 => x"3306c500",
        3410 => x"6316c500",
        3411 => x"13050000",
        3412 => x"67800000",
        3413 => x"83470500",
        3414 => x"e38cb7fe",
        3415 => x"13051500",
        3416 => x"6ff09ffe",
        3417 => x"130101ff",
        3418 => x"23248100",
        3419 => x"23229100",
        3420 => x"13040500",
        3421 => x"13850500",
        3422 => x"93050600",
        3423 => x"23261100",
        3424 => x"23a20188",
        3425 => x"efd0dfe2",
        3426 => x"9307f0ff",
        3427 => x"6318f500",
        3428 => x"83a74188",
        3429 => x"63840700",
        3430 => x"2320f400",
        3431 => x"8320c100",
        3432 => x"03248100",
        3433 => x"83244100",
        3434 => x"13010101",
        3435 => x"67800000",
        3436 => x"130101ff",
        3437 => x"23248100",
        3438 => x"23229100",
        3439 => x"13040500",
        3440 => x"13850500",
        3441 => x"23261100",
        3442 => x"23a20188",
        3443 => x"efe00f86",
        3444 => x"9307f0ff",
        3445 => x"6318f500",
        3446 => x"83a74188",
        3447 => x"63840700",
        3448 => x"2320f400",
        3449 => x"8320c100",
        3450 => x"03248100",
        3451 => x"83244100",
        3452 => x"13010101",
        3453 => x"67800000",
        3454 => x"130101fe",
        3455 => x"232c8100",
        3456 => x"232e1100",
        3457 => x"232a9100",
        3458 => x"23282101",
        3459 => x"23263101",
        3460 => x"23244101",
        3461 => x"13040600",
        3462 => x"63940502",
        3463 => x"03248101",
        3464 => x"8320c101",
        3465 => x"83244101",
        3466 => x"03290101",
        3467 => x"8329c100",
        3468 => x"032a8100",
        3469 => x"93050600",
        3470 => x"13010102",
        3471 => x"6fe05fec",
        3472 => x"63180602",
        3473 => x"efe01fd4",
        3474 => x"93040000",
        3475 => x"8320c101",
        3476 => x"03248101",
        3477 => x"03290101",
        3478 => x"8329c100",
        3479 => x"032a8100",
        3480 => x"13850400",
        3481 => x"83244101",
        3482 => x"13010102",
        3483 => x"67800000",
        3484 => x"130a0500",
        3485 => x"93840500",
        3486 => x"ef008005",
        3487 => x"13090500",
        3488 => x"63668500",
        3489 => x"93571500",
        3490 => x"e3e287fc",
        3491 => x"93050400",
        3492 => x"13050a00",
        3493 => x"efe0dfe6",
        3494 => x"93090500",
        3495 => x"63160500",
        3496 => x"93840900",
        3497 => x"6ff09ffa",
        3498 => x"13060400",
        3499 => x"63748900",
        3500 => x"13060900",
        3501 => x"93850400",
        3502 => x"13850900",
        3503 => x"efd01fc9",
        3504 => x"93850400",
        3505 => x"13050a00",
        3506 => x"efe0dfcb",
        3507 => x"6ff05ffd",
        3508 => x"83a7c5ff",
        3509 => x"1385c7ff",
        3510 => x"63d80700",
        3511 => x"b385a500",
        3512 => x"83a70500",
        3513 => x"3305f500",
        3514 => x"67800000",
        3515 => x"10000000",
        3516 => x"00000000",
        3517 => x"037a5200",
        3518 => x"017c0101",
        3519 => x"1b0d0200",
        3520 => x"10000000",
        3521 => x"18000000",
        3522 => x"9ccfffff",
        3523 => x"78040000",
        3524 => x"00000000",
        3525 => x"10000000",
        3526 => x"00000000",
        3527 => x"037a5200",
        3528 => x"017c0101",
        3529 => x"1b0d0200",
        3530 => x"10000000",
        3531 => x"18000000",
        3532 => x"ecd3ffff",
        3533 => x"30040000",
        3534 => x"00000000",
        3535 => x"10000000",
        3536 => x"00000000",
        3537 => x"037a5200",
        3538 => x"017c0101",
        3539 => x"1b0d0200",
        3540 => x"10000000",
        3541 => x"18000000",
        3542 => x"f4d7ffff",
        3543 => x"e4030000",
        3544 => x"00000000",
        3545 => x"30313233",
        3546 => x"34353637",
        3547 => x"38396162",
        3548 => x"63646566",
        3549 => x"00000000",
        3550 => x"64040000",
        3551 => x"9c030000",
        3552 => x"9c030000",
        3553 => x"9c030000",
        3554 => x"9c030000",
        3555 => x"9c030000",
        3556 => x"9c030000",
        3557 => x"9c030000",
        3558 => x"9c030000",
        3559 => x"70040000",
        3560 => x"7c040000",
        3561 => x"88040000",
        3562 => x"94040000",
        3563 => x"a0040000",
        3564 => x"58040000",
        3565 => x"9c030000",
        3566 => x"9c030000",
        3567 => x"9c030000",
        3568 => x"ac040000",
        3569 => x"9c030000",
        3570 => x"9c030000",
        3571 => x"9c030000",
        3572 => x"9c030000",
        3573 => x"9c030000",
        3574 => x"9c030000",
        3575 => x"9c030000",
        3576 => x"bc040000",
        3577 => x"50050000",
        3578 => x"68050000",
        3579 => x"98050000",
        3580 => x"18050000",
        3581 => x"18050000",
        3582 => x"18050000",
        3583 => x"18050000",
        3584 => x"18050000",
        3585 => x"18050000",
        3586 => x"80050000",
        3587 => x"18050000",
        3588 => x"18050000",
        3589 => x"18050000",
        3590 => x"18050000",
        3591 => x"30050000",
        3592 => x"30050000",
        3593 => x"50050000",
        3594 => x"18050000",
        3595 => x"18050000",
        3596 => x"18050000",
        3597 => x"18050000",
        3598 => x"44050000",
        3599 => x"b0050000",
        3600 => x"d8050000",
        3601 => x"18050000",
        3602 => x"18050000",
        3603 => x"18050000",
        3604 => x"18050000",
        3605 => x"18050000",
        3606 => x"18050000",
        3607 => x"18050000",
        3608 => x"18050000",
        3609 => x"18050000",
        3610 => x"18050000",
        3611 => x"18050000",
        3612 => x"18050000",
        3613 => x"18050000",
        3614 => x"18050000",
        3615 => x"30050000",
        3616 => x"30050000",
        3617 => x"18050000",
        3618 => x"18050000",
        3619 => x"18050000",
        3620 => x"18050000",
        3621 => x"18050000",
        3622 => x"18050000",
        3623 => x"18050000",
        3624 => x"18050000",
        3625 => x"18050000",
        3626 => x"18050000",
        3627 => x"18050000",
        3628 => x"18050000",
        3629 => x"44050000",
        3630 => x"00010202",
        3631 => x"03030303",
        3632 => x"04040404",
        3633 => x"04040404",
        3634 => x"05050505",
        3635 => x"05050505",
        3636 => x"05050505",
        3637 => x"05050505",
        3638 => x"06060606",
        3639 => x"06060606",
        3640 => x"06060606",
        3641 => x"06060606",
        3642 => x"06060606",
        3643 => x"06060606",
        3644 => x"06060606",
        3645 => x"06060606",
        3646 => x"07070707",
        3647 => x"07070707",
        3648 => x"07070707",
        3649 => x"07070707",
        3650 => x"07070707",
        3651 => x"07070707",
        3652 => x"07070707",
        3653 => x"07070707",
        3654 => x"07070707",
        3655 => x"07070707",
        3656 => x"07070707",
        3657 => x"07070707",
        3658 => x"07070707",
        3659 => x"07070707",
        3660 => x"07070707",
        3661 => x"07070707",
        3662 => x"08080808",
        3663 => x"08080808",
        3664 => x"08080808",
        3665 => x"08080808",
        3666 => x"08080808",
        3667 => x"08080808",
        3668 => x"08080808",
        3669 => x"08080808",
        3670 => x"08080808",
        3671 => x"08080808",
        3672 => x"08080808",
        3673 => x"08080808",
        3674 => x"08080808",
        3675 => x"08080808",
        3676 => x"08080808",
        3677 => x"08080808",
        3678 => x"08080808",
        3679 => x"08080808",
        3680 => x"08080808",
        3681 => x"08080808",
        3682 => x"08080808",
        3683 => x"08080808",
        3684 => x"08080808",
        3685 => x"08080808",
        3686 => x"08080808",
        3687 => x"08080808",
        3688 => x"08080808",
        3689 => x"08080808",
        3690 => x"08080808",
        3691 => x"08080808",
        3692 => x"08080808",
        3693 => x"08080808",
        3694 => x"0d0a4542",
        3695 => x"5245414b",
        3696 => x"21206d65",
        3697 => x"7063203d",
        3698 => x"20000000",
        3699 => x"20696e73",
        3700 => x"6e203d20",
        3701 => x"00000000",
        3702 => x"0d0a0d0a",
        3703 => x"44697370",
        3704 => x"6c617969",
        3705 => x"6e672074",
        3706 => x"68652074",
        3707 => x"696d6520",
        3708 => x"70617373",
        3709 => x"65642073",
        3710 => x"696e6365",
        3711 => x"20726573",
        3712 => x"65740d0a",
        3713 => x"0d0a0000",
        3714 => x"2530356c",
        3715 => x"643a2530",
        3716 => x"366c6420",
        3717 => x"20202530",
        3718 => x"326c643a",
        3719 => x"2530326c",
        3720 => x"643a2530",
        3721 => x"326c640d",
        3722 => x"00000000",
        3723 => x"696e7465",
        3724 => x"72727570",
        3725 => x"745f6469",
        3726 => x"72656374",
        3727 => x"00000000",
        3728 => x"54485541",
        3729 => x"53205249",
        3730 => x"53432d56",
        3731 => x"20525633",
        3732 => x"32494d20",
        3733 => x"62617265",
        3734 => x"206d6574",
        3735 => x"616c2070",
        3736 => x"726f6365",
        3737 => x"73736f72",
        3738 => x"00000000",
        3739 => x"54686520",
        3740 => x"48616775",
        3741 => x"6520556e",
        3742 => x"69766572",
        3743 => x"73697479",
        3744 => x"206f6620",
        3745 => x"4170706c",
        3746 => x"69656420",
        3747 => x"53636965",
        3748 => x"6e636573",
        3749 => x"00000000",
        3750 => x"44657061",
        3751 => x"72746d65",
        3752 => x"6e74206f",
        3753 => x"6620456c",
        3754 => x"65637472",
        3755 => x"6963616c",
        3756 => x"20456e67",
        3757 => x"696e6565",
        3758 => x"72696e67",
        3759 => x"00000000",
        3760 => x"4a2e452e",
        3761 => x"4a2e206f",
        3762 => x"70206465",
        3763 => x"6e204272",
        3764 => x"6f757700",
        3765 => x"232d302b",
        3766 => x"20000000",
        3767 => x"686c4c00",
        3768 => x"65666745",
        3769 => x"46470000",
        3770 => x"30313233",
        3771 => x"34353637",
        3772 => x"38394142",
        3773 => x"43444546",
        3774 => x"00000000",
        3775 => x"30313233",
        3776 => x"34353637",
        3777 => x"38396162",
        3778 => x"63646566",
        3779 => x"00000000",
        3780 => x"cc2f0000",
        3781 => x"ec2f0000",
        3782 => x"982f0000",
        3783 => x"982f0000",
        3784 => x"982f0000",
        3785 => x"982f0000",
        3786 => x"ec2f0000",
        3787 => x"982f0000",
        3788 => x"982f0000",
        3789 => x"982f0000",
        3790 => x"982f0000",
        3791 => x"d8310000",
        3792 => x"44300000",
        3793 => x"50310000",
        3794 => x"982f0000",
        3795 => x"982f0000",
        3796 => x"20320000",
        3797 => x"982f0000",
        3798 => x"44300000",
        3799 => x"982f0000",
        3800 => x"982f0000",
        3801 => x"5c310000",
        3802 => x"2c3a0000",
        3803 => x"403a0000",
        3804 => x"6c3a0000",
        3805 => x"983a0000",
        3806 => x"c03a0000",
        3807 => x"00000000",
        3808 => x"00000000",
        3809 => x"03000000",
        3810 => x"90000020",
        3811 => x"00000000",
        3812 => x"90000020",
        3813 => x"f8000020",
        3814 => x"60010020",
        3815 => x"00000000",
        3816 => x"00000000",
        3817 => x"00000000",
        3818 => x"00000000",
        3819 => x"00000000",
        3820 => x"00000000",
        3821 => x"00000000",
        3822 => x"00000000",
        3823 => x"00000000",
        3824 => x"00000000",
        3825 => x"00000000",
        3826 => x"00000000",
        3827 => x"00000000",
        3828 => x"00000000",
        3829 => x"00000000",
        3830 => x"78000020",
        3831 => x"24000020"
            );
end package rom_image;
