-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Tue Dec 17 09:18:29 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382c22e",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"13060500",
           9 => x"93874187",
          10 => x"637cf600",
          11 => x"b7450000",
          12 => x"3386c740",
          13 => x"13050500",
          14 => x"9385c5c4",
          15 => x"ef10003e",
          16 => x"13864187",
          17 => x"9387019c",
          18 => x"637af600",
          19 => x"3386c740",
          20 => x"13854187",
          21 => x"93050000",
          22 => x"ef10803a",
          23 => x"ef208011",
          24 => x"b7050020",
          25 => x"93850500",
          26 => x"13060000",
          27 => x"13055000",
          28 => x"ef10c04b",
          29 => x"ef109008",
          30 => x"6f104040",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef108044",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"b7470000",
          40 => x"232c4101",
          41 => x"130a0500",
          42 => x"138507a6",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"37390000",
          50 => x"ef104042",
          51 => x"13044100",
          52 => x"93070400",
          53 => x"9309c1ff",
          54 => x"1309497e",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef10c03e",
          65 => x"37450000",
          66 => x"130545a7",
          67 => x"ef10003e",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef10803b",
          78 => x"37450000",
          79 => x"130505a8",
          80 => x"ef10c03a",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74760",
          91 => x"93860700",
          92 => x"1377f7fe",
          93 => x"23a2e760",
          94 => x"83a74700",
          95 => x"93c71700",
          96 => x"23a2f600",
          97 => x"67800000",
          98 => x"370700f0",
          99 => x"83274700",
         100 => x"93e70720",
         101 => x"2322f700",
         102 => x"6f000000",
         103 => x"b71700f0",
         104 => x"93850700",
         105 => x"938505a0",
         106 => x"938747a0",
         107 => x"83a60700",
         108 => x"03a60500",
         109 => x"03a70700",
         110 => x"e31ad7fe",
         111 => x"b7870100",
         112 => x"b71600f0",
         113 => x"1305f0ff",
         114 => x"9387076a",
         115 => x"23a6a6a0",
         116 => x"b307f600",
         117 => x"23a4a6a0",
         118 => x"33b6c700",
         119 => x"23a4f6a0",
         120 => x"3306e600",
         121 => x"23a6c6a0",
         122 => x"370700f0",
         123 => x"83274700",
         124 => x"93c72700",
         125 => x"2322f700",
         126 => x"67800000",
         127 => x"b70700f0",
         128 => x"03a74710",
         129 => x"b70600f0",
         130 => x"93870710",
         131 => x"13778700",
         132 => x"630a0700",
         133 => x"03a74600",
         134 => x"13478700",
         135 => x"23a2e600",
         136 => x"83a78700",
         137 => x"67800000",
         138 => x"b70700f0",
         139 => x"03a74770",
         140 => x"93860700",
         141 => x"1377f7f0",
         142 => x"23a2e770",
         143 => x"83a74700",
         144 => x"93c74700",
         145 => x"23a2f600",
         146 => x"67800000",
         147 => x"b70700f0",
         148 => x"03a74740",
         149 => x"93860700",
         150 => x"137777ff",
         151 => x"23a2e740",
         152 => x"83a74700",
         153 => x"93c70701",
         154 => x"23a2f600",
         155 => x"67800000",
         156 => x"b70700f0",
         157 => x"03a74720",
         158 => x"93860700",
         159 => x"137777ff",
         160 => x"23a2e720",
         161 => x"83a74700",
         162 => x"93c70702",
         163 => x"23a2f600",
         164 => x"67800000",
         165 => x"b70700f0",
         166 => x"03a74730",
         167 => x"93860700",
         168 => x"137777ff",
         169 => x"23a2e730",
         170 => x"83a74700",
         171 => x"93c70708",
         172 => x"23a2f600",
         173 => x"67800000",
         174 => x"b70700f0",
         175 => x"23ae0700",
         176 => x"03a74700",
         177 => x"13470704",
         178 => x"23a2e700",
         179 => x"67800000",
         180 => x"b71700f0",
         181 => x"23a00790",
         182 => x"370700f0",
         183 => x"83274700",
         184 => x"93c70710",
         185 => x"2322f700",
         186 => x"67800000",
         187 => x"6f000000",
         188 => x"13050000",
         189 => x"67800000",
         190 => x"13050000",
         191 => x"67800000",
         192 => x"130101f7",
         193 => x"23221100",
         194 => x"23242100",
         195 => x"23263100",
         196 => x"23284100",
         197 => x"232a5100",
         198 => x"232c6100",
         199 => x"232e7100",
         200 => x"23208102",
         201 => x"23229102",
         202 => x"2324a102",
         203 => x"2326b102",
         204 => x"2328c102",
         205 => x"232ad102",
         206 => x"232ce102",
         207 => x"232ef102",
         208 => x"23200105",
         209 => x"23221105",
         210 => x"23242105",
         211 => x"23263105",
         212 => x"23284105",
         213 => x"232a5105",
         214 => x"232c6105",
         215 => x"232e7105",
         216 => x"23208107",
         217 => x"23229107",
         218 => x"2324a107",
         219 => x"2326b107",
         220 => x"2328c107",
         221 => x"232ad107",
         222 => x"232ce107",
         223 => x"232ef107",
         224 => x"f3222034",
         225 => x"23205108",
         226 => x"f3221034",
         227 => x"23225108",
         228 => x"83a20200",
         229 => x"23245108",
         230 => x"f3223034",
         231 => x"23265108",
         232 => x"f3272034",
         233 => x"1307b000",
         234 => x"6374f70c",
         235 => x"37070080",
         236 => x"1307d7ff",
         237 => x"b387e700",
         238 => x"13078001",
         239 => x"636ef700",
         240 => x"37370000",
         241 => x"93972700",
         242 => x"1307877f",
         243 => x"b387e700",
         244 => x"83a70700",
         245 => x"67800700",
         246 => x"03258102",
         247 => x"83220108",
         248 => x"63c80200",
         249 => x"f3221034",
         250 => x"93824200",
         251 => x"73901234",
         252 => x"832fc107",
         253 => x"032f8107",
         254 => x"832e4107",
         255 => x"032e0107",
         256 => x"832dc106",
         257 => x"032d8106",
         258 => x"832c4106",
         259 => x"032c0106",
         260 => x"832bc105",
         261 => x"032b8105",
         262 => x"832a4105",
         263 => x"032a0105",
         264 => x"8329c104",
         265 => x"03298104",
         266 => x"83284104",
         267 => x"03280104",
         268 => x"8327c103",
         269 => x"03278103",
         270 => x"83264103",
         271 => x"03260103",
         272 => x"8325c102",
         273 => x"83244102",
         274 => x"03240102",
         275 => x"8323c101",
         276 => x"03238101",
         277 => x"83224101",
         278 => x"03220101",
         279 => x"8321c100",
         280 => x"03218100",
         281 => x"83204100",
         282 => x"13010109",
         283 => x"73002030",
         284 => x"93061000",
         285 => x"e3f2f6f6",
         286 => x"e360f7f6",
         287 => x"37470000",
         288 => x"93972700",
         289 => x"1307c785",
         290 => x"b387e700",
         291 => x"83a70700",
         292 => x"67800700",
         293 => x"eff09fdb",
         294 => x"03258102",
         295 => x"6ff01ff4",
         296 => x"eff01fe3",
         297 => x"03258102",
         298 => x"6ff05ff3",
         299 => x"eff01fcf",
         300 => x"03258102",
         301 => x"6ff09ff2",
         302 => x"eff01fe0",
         303 => x"03258102",
         304 => x"6ff0dff1",
         305 => x"eff01fca",
         306 => x"03258102",
         307 => x"6ff01ff1",
         308 => x"eff09fd5",
         309 => x"03258102",
         310 => x"6ff05ff0",
         311 => x"eff01fd2",
         312 => x"03258102",
         313 => x"6ff09fef",
         314 => x"eff0dfda",
         315 => x"03258102",
         316 => x"6ff0dfee",
         317 => x"eff0dfd7",
         318 => x"03258102",
         319 => x"6ff01fee",
         320 => x"13050100",
         321 => x"eff05fb9",
         322 => x"03258102",
         323 => x"6ff01fed",
         324 => x"9307600d",
         325 => x"6380f81c",
         326 => x"63cc1703",
         327 => x"9307d005",
         328 => x"63c21715",
         329 => x"93078003",
         330 => x"63da1705",
         331 => x"938878fc",
         332 => x"93074002",
         333 => x"63e41705",
         334 => x"b7470000",
         335 => x"9387c788",
         336 => x"93982800",
         337 => x"b388f800",
         338 => x"83a70800",
         339 => x"67800700",
         340 => x"93073019",
         341 => x"6388f818",
         342 => x"938808c0",
         343 => x"9307f000",
         344 => x"63ee1701",
         345 => x"b7470000",
         346 => x"93870792",
         347 => x"93982800",
         348 => x"b388f800",
         349 => x"83a70800",
         350 => x"67800700",
         351 => x"ef10103f",
         352 => x"93078005",
         353 => x"2320f500",
         354 => x"9307f0ff",
         355 => x"13850700",
         356 => x"6ff0dfe4",
         357 => x"b7270000",
         358 => x"23a2f500",
         359 => x"93070000",
         360 => x"13850700",
         361 => x"6ff09fe3",
         362 => x"ef10503c",
         363 => x"93079000",
         364 => x"2320f500",
         365 => x"9307f0ff",
         366 => x"13850700",
         367 => x"6ff01fe2",
         368 => x"ef10d03a",
         369 => x"9307d000",
         370 => x"2320f500",
         371 => x"9307f0ff",
         372 => x"13850700",
         373 => x"6ff09fe0",
         374 => x"ef105039",
         375 => x"93072000",
         376 => x"2320f500",
         377 => x"9307f0ff",
         378 => x"13850700",
         379 => x"6ff01fdf",
         380 => x"ef10d037",
         381 => x"9307f001",
         382 => x"2320f500",
         383 => x"9307f0ff",
         384 => x"13850700",
         385 => x"6ff09fdd",
         386 => x"93070000",
         387 => x"13850700",
         388 => x"6ff0dfdc",
         389 => x"13090600",
         390 => x"13840500",
         391 => x"635cc000",
         392 => x"b384c500",
         393 => x"03450400",
         394 => x"13041400",
         395 => x"eff01fa5",
         396 => x"e39a84fe",
         397 => x"13050900",
         398 => x"6ff05fda",
         399 => x"13090600",
         400 => x"13840500",
         401 => x"e358c0fe",
         402 => x"b384c500",
         403 => x"eff0dfa2",
         404 => x"2300a400",
         405 => x"13041400",
         406 => x"e39a84fe",
         407 => x"13050900",
         408 => x"6ff0dfd7",
         409 => x"9307900a",
         410 => x"e39af8f0",
         411 => x"13090000",
         412 => x"93040500",
         413 => x"13040900",
         414 => x"93090900",
         415 => x"93070900",
         416 => x"732410c8",
         417 => x"f32910c0",
         418 => x"f32710c8",
         419 => x"e31af4fe",
         420 => x"37460f00",
         421 => x"13060624",
         422 => x"93060000",
         423 => x"13850900",
         424 => x"93050400",
         425 => x"ef00d017",
         426 => x"37460f00",
         427 => x"23a4a400",
         428 => x"93050400",
         429 => x"13850900",
         430 => x"13060624",
         431 => x"93060000",
         432 => x"ef004053",
         433 => x"23a0a400",
         434 => x"23a2b400",
         435 => x"13050900",
         436 => x"6ff0dfd0",
         437 => x"63100508",
         438 => x"1385019c",
         439 => x"13050500",
         440 => x"6ff0dfcf",
         441 => x"13090000",
         442 => x"93840500",
         443 => x"13040900",
         444 => x"93090900",
         445 => x"93070900",
         446 => x"732410c8",
         447 => x"f32910c0",
         448 => x"f32710c8",
         449 => x"e31af4fe",
         450 => x"37460f00",
         451 => x"13060624",
         452 => x"93060000",
         453 => x"13850900",
         454 => x"93050400",
         455 => x"ef005010",
         456 => x"9307803e",
         457 => x"b307f502",
         458 => x"37460f00",
         459 => x"93050400",
         460 => x"13850900",
         461 => x"13060624",
         462 => x"93060000",
         463 => x"23a4f400",
         464 => x"ef00404b",
         465 => x"23a0a400",
         466 => x"23a2b400",
         467 => x"13050900",
         468 => x"6ff0dfc8",
         469 => x"b7870020",
         470 => x"93870700",
         471 => x"13070040",
         472 => x"b387e740",
         473 => x"e36cf5f6",
         474 => x"ef105020",
         475 => x"9307c000",
         476 => x"2320f500",
         477 => x"1305f0ff",
         478 => x"13050500",
         479 => x"6ff01fc6",
         480 => x"13030500",
         481 => x"138e0500",
         482 => x"93080000",
         483 => x"63dc0500",
         484 => x"b337a000",
         485 => x"3307b040",
         486 => x"330ef740",
         487 => x"3303a040",
         488 => x"9308f0ff",
         489 => x"63dc0600",
         490 => x"b337c000",
         491 => x"b306d040",
         492 => x"93c8f8ff",
         493 => x"b386f640",
         494 => x"3306c040",
         495 => x"13070600",
         496 => x"13080300",
         497 => x"93070e00",
         498 => x"639c0628",
         499 => x"b7450000",
         500 => x"93850596",
         501 => x"6376ce0e",
         502 => x"b7060100",
         503 => x"6378d60c",
         504 => x"93360610",
         505 => x"93b61600",
         506 => x"93963600",
         507 => x"3355d600",
         508 => x"b385a500",
         509 => x"83c50500",
         510 => x"13050002",
         511 => x"b386d500",
         512 => x"b305d540",
         513 => x"630cd500",
         514 => x"b317be00",
         515 => x"b356d300",
         516 => x"3317b600",
         517 => x"b3e7f600",
         518 => x"3318b300",
         519 => x"93550701",
         520 => x"33deb702",
         521 => x"13160701",
         522 => x"13560601",
         523 => x"b3f7b702",
         524 => x"13050e00",
         525 => x"3303c603",
         526 => x"93960701",
         527 => x"93570801",
         528 => x"b3e7d700",
         529 => x"63fe6700",
         530 => x"b307f700",
         531 => x"1305feff",
         532 => x"63e8e700",
         533 => x"63f66700",
         534 => x"1305eeff",
         535 => x"b387e700",
         536 => x"b3876740",
         537 => x"33d3b702",
         538 => x"13180801",
         539 => x"13580801",
         540 => x"b3f7b702",
         541 => x"b3066602",
         542 => x"93970701",
         543 => x"3368f800",
         544 => x"93070300",
         545 => x"637cd800",
         546 => x"33080701",
         547 => x"9307f3ff",
         548 => x"6366e800",
         549 => x"6374d800",
         550 => x"9307e3ff",
         551 => x"13150501",
         552 => x"3365f500",
         553 => x"93050000",
         554 => x"6f00000e",
         555 => x"37050001",
         556 => x"93068001",
         557 => x"e37ca6f2",
         558 => x"93060001",
         559 => x"6ff01ff3",
         560 => x"93060000",
         561 => x"630c0600",
         562 => x"b7070100",
         563 => x"637af60c",
         564 => x"93360610",
         565 => x"93b61600",
         566 => x"93963600",
         567 => x"b357d600",
         568 => x"b385f500",
         569 => x"83c70500",
         570 => x"b387d700",
         571 => x"93060002",
         572 => x"b385f640",
         573 => x"6390f60c",
         574 => x"b307ce40",
         575 => x"93051000",
         576 => x"13530701",
         577 => x"b3de6702",
         578 => x"13160701",
         579 => x"13560601",
         580 => x"93560801",
         581 => x"b3f76702",
         582 => x"13850e00",
         583 => x"330ed603",
         584 => x"93970701",
         585 => x"b3e7f600",
         586 => x"63fec701",
         587 => x"b307f700",
         588 => x"1385feff",
         589 => x"63e8e700",
         590 => x"63f6c701",
         591 => x"1385eeff",
         592 => x"b387e700",
         593 => x"b387c741",
         594 => x"33de6702",
         595 => x"13180801",
         596 => x"13580801",
         597 => x"b3f76702",
         598 => x"b306c603",
         599 => x"93970701",
         600 => x"3368f800",
         601 => x"93070e00",
         602 => x"637cd800",
         603 => x"33080701",
         604 => x"9307feff",
         605 => x"6366e800",
         606 => x"6374d800",
         607 => x"9307eeff",
         608 => x"13150501",
         609 => x"3365f500",
         610 => x"638a0800",
         611 => x"b337a000",
         612 => x"b305b040",
         613 => x"b385f540",
         614 => x"3305a040",
         615 => x"67800000",
         616 => x"b7070001",
         617 => x"93068001",
         618 => x"e37af6f2",
         619 => x"93060001",
         620 => x"6ff0dff2",
         621 => x"3317b600",
         622 => x"b356fe00",
         623 => x"13550701",
         624 => x"331ebe00",
         625 => x"b357f300",
         626 => x"b3e7c701",
         627 => x"33dea602",
         628 => x"13160701",
         629 => x"13560601",
         630 => x"3318b300",
         631 => x"b3f6a602",
         632 => x"3303c603",
         633 => x"93950601",
         634 => x"93d60701",
         635 => x"b3e6b600",
         636 => x"93050e00",
         637 => x"63fe6600",
         638 => x"b306d700",
         639 => x"9305feff",
         640 => x"63e8e600",
         641 => x"63f66600",
         642 => x"9305eeff",
         643 => x"b386e600",
         644 => x"b3866640",
         645 => x"33d3a602",
         646 => x"93970701",
         647 => x"93d70701",
         648 => x"b3f6a602",
         649 => x"33066602",
         650 => x"93960601",
         651 => x"b3e7d700",
         652 => x"93060300",
         653 => x"63fec700",
         654 => x"b307f700",
         655 => x"9306f3ff",
         656 => x"63e8e700",
         657 => x"63f6c700",
         658 => x"9306e3ff",
         659 => x"b387e700",
         660 => x"93950501",
         661 => x"b387c740",
         662 => x"b3e5d500",
         663 => x"6ff05fea",
         664 => x"6364de18",
         665 => x"b7070100",
         666 => x"63f4f604",
         667 => x"13b70610",
         668 => x"13371700",
         669 => x"13173700",
         670 => x"b7470000",
         671 => x"b3d5e600",
         672 => x"93870796",
         673 => x"b387b700",
         674 => x"83c70700",
         675 => x"b387e700",
         676 => x"13070002",
         677 => x"b305f740",
         678 => x"6316f702",
         679 => x"13051000",
         680 => x"e3e4c6ef",
         681 => x"3335c300",
         682 => x"13351500",
         683 => x"6ff0dfed",
         684 => x"b7070001",
         685 => x"13078001",
         686 => x"e3f0f6fc",
         687 => x"13070001",
         688 => x"6ff09ffb",
         689 => x"3358f600",
         690 => x"b396b600",
         691 => x"3368d800",
         692 => x"3355fe00",
         693 => x"3317be00",
         694 => x"135e0801",
         695 => x"335fc503",
         696 => x"93160801",
         697 => x"93d60601",
         698 => x"b357f300",
         699 => x"b3e7e700",
         700 => x"13d70701",
         701 => x"3316b600",
         702 => x"3375c503",
         703 => x"b38ee603",
         704 => x"13150501",
         705 => x"3367a700",
         706 => x"13050f00",
         707 => x"637ed701",
         708 => x"3307e800",
         709 => x"1305ffff",
         710 => x"63680701",
         711 => x"6376d701",
         712 => x"1305efff",
         713 => x"33070701",
         714 => x"3307d741",
         715 => x"b35ec703",
         716 => x"93970701",
         717 => x"93d70701",
         718 => x"3377c703",
         719 => x"b386d603",
         720 => x"13170701",
         721 => x"b3e7e700",
         722 => x"13870e00",
         723 => x"63fed700",
         724 => x"b307f800",
         725 => x"1387feff",
         726 => x"63e80701",
         727 => x"63f6d700",
         728 => x"1387eeff",
         729 => x"b3870701",
         730 => x"13150501",
         731 => x"3365e500",
         732 => x"131e0601",
         733 => x"13170701",
         734 => x"13570701",
         735 => x"13580501",
         736 => x"135e0e01",
         737 => x"13560601",
         738 => x"b30ec703",
         739 => x"b387d740",
         740 => x"330ec803",
         741 => x"93d60e01",
         742 => x"3307c702",
         743 => x"3307c701",
         744 => x"3387e600",
         745 => x"3308c802",
         746 => x"6376c701",
         747 => x"b7060100",
         748 => x"3308d800",
         749 => x"93560701",
         750 => x"b3860601",
         751 => x"63e2d702",
         752 => x"e392d7ce",
         753 => x"939e0e01",
         754 => x"13170701",
         755 => x"93de0e01",
         756 => x"3313b300",
         757 => x"3307d701",
         758 => x"93050000",
         759 => x"e376e3da",
         760 => x"1305f5ff",
         761 => x"6ff01fcc",
         762 => x"93050000",
         763 => x"13050000",
         764 => x"6ff09fd9",
         765 => x"93080500",
         766 => x"13830500",
         767 => x"13070600",
         768 => x"13080500",
         769 => x"93870500",
         770 => x"63920628",
         771 => x"b7450000",
         772 => x"93850596",
         773 => x"6376c30e",
         774 => x"b7060100",
         775 => x"6378d60c",
         776 => x"93360610",
         777 => x"93b61600",
         778 => x"93963600",
         779 => x"3355d600",
         780 => x"b385a500",
         781 => x"83c50500",
         782 => x"13050002",
         783 => x"b386d500",
         784 => x"b305d540",
         785 => x"630cd500",
         786 => x"b317b300",
         787 => x"b3d6d800",
         788 => x"3317b600",
         789 => x"b3e7f600",
         790 => x"3398b800",
         791 => x"93550701",
         792 => x"33d3b702",
         793 => x"13160701",
         794 => x"13560601",
         795 => x"b3f7b702",
         796 => x"13050300",
         797 => x"b3086602",
         798 => x"93960701",
         799 => x"93570801",
         800 => x"b3e7d700",
         801 => x"63fe1701",
         802 => x"b307f700",
         803 => x"1305f3ff",
         804 => x"63e8e700",
         805 => x"63f61701",
         806 => x"1305e3ff",
         807 => x"b387e700",
         808 => x"b3871741",
         809 => x"b3d8b702",
         810 => x"13180801",
         811 => x"13580801",
         812 => x"b3f7b702",
         813 => x"b3061603",
         814 => x"93970701",
         815 => x"3368f800",
         816 => x"93870800",
         817 => x"637cd800",
         818 => x"33080701",
         819 => x"9387f8ff",
         820 => x"6366e800",
         821 => x"6374d800",
         822 => x"9387e8ff",
         823 => x"13150501",
         824 => x"3365f500",
         825 => x"93050000",
         826 => x"67800000",
         827 => x"37050001",
         828 => x"93068001",
         829 => x"e37ca6f2",
         830 => x"93060001",
         831 => x"6ff01ff3",
         832 => x"93060000",
         833 => x"630c0600",
         834 => x"b7070100",
         835 => x"6370f60c",
         836 => x"93360610",
         837 => x"93b61600",
         838 => x"93963600",
         839 => x"b357d600",
         840 => x"b385f500",
         841 => x"83c70500",
         842 => x"b387d700",
         843 => x"93060002",
         844 => x"b385f640",
         845 => x"6396f60a",
         846 => x"b307c340",
         847 => x"93051000",
         848 => x"93580701",
         849 => x"33de1703",
         850 => x"13160701",
         851 => x"13560601",
         852 => x"93560801",
         853 => x"b3f71703",
         854 => x"13050e00",
         855 => x"3303c603",
         856 => x"93970701",
         857 => x"b3e7f600",
         858 => x"63fe6700",
         859 => x"b307f700",
         860 => x"1305feff",
         861 => x"63e8e700",
         862 => x"63f66700",
         863 => x"1305eeff",
         864 => x"b387e700",
         865 => x"b3876740",
         866 => x"33d31703",
         867 => x"13180801",
         868 => x"13580801",
         869 => x"b3f71703",
         870 => x"b3066602",
         871 => x"93970701",
         872 => x"3368f800",
         873 => x"93070300",
         874 => x"637cd800",
         875 => x"33080701",
         876 => x"9307f3ff",
         877 => x"6366e800",
         878 => x"6374d800",
         879 => x"9307e3ff",
         880 => x"13150501",
         881 => x"3365f500",
         882 => x"67800000",
         883 => x"b7070001",
         884 => x"93068001",
         885 => x"e374f6f4",
         886 => x"93060001",
         887 => x"6ff01ff4",
         888 => x"3317b600",
         889 => x"b356f300",
         890 => x"13550701",
         891 => x"3313b300",
         892 => x"b3d7f800",
         893 => x"b3e76700",
         894 => x"33d3a602",
         895 => x"13160701",
         896 => x"13560601",
         897 => x"3398b800",
         898 => x"b3f6a602",
         899 => x"b3086602",
         900 => x"93950601",
         901 => x"93d60701",
         902 => x"b3e6b600",
         903 => x"93050300",
         904 => x"63fe1601",
         905 => x"b306d700",
         906 => x"9305f3ff",
         907 => x"63e8e600",
         908 => x"63f61601",
         909 => x"9305e3ff",
         910 => x"b386e600",
         911 => x"b3861641",
         912 => x"b3d8a602",
         913 => x"93970701",
         914 => x"93d70701",
         915 => x"b3f6a602",
         916 => x"33061603",
         917 => x"93960601",
         918 => x"b3e7d700",
         919 => x"93860800",
         920 => x"63fec700",
         921 => x"b307f700",
         922 => x"9386f8ff",
         923 => x"63e8e700",
         924 => x"63f6c700",
         925 => x"9386e8ff",
         926 => x"b387e700",
         927 => x"93950501",
         928 => x"b387c740",
         929 => x"b3e5d500",
         930 => x"6ff09feb",
         931 => x"63e4d518",
         932 => x"b7070100",
         933 => x"63f4f604",
         934 => x"93b70610",
         935 => x"93b71700",
         936 => x"93973700",
         937 => x"37470000",
         938 => x"b3d5f600",
         939 => x"13070796",
         940 => x"3307b700",
         941 => x"03470700",
         942 => x"3307f700",
         943 => x"93070002",
         944 => x"b385e740",
         945 => x"6396e702",
         946 => x"13051000",
         947 => x"e3ee66e0",
         948 => x"33b5c800",
         949 => x"13351500",
         950 => x"67800000",
         951 => x"37070001",
         952 => x"93078001",
         953 => x"e3f0e6fc",
         954 => x"93070001",
         955 => x"6ff09ffb",
         956 => x"3355e600",
         957 => x"b396b600",
         958 => x"b357e300",
         959 => x"3365d500",
         960 => x"3313b300",
         961 => x"33d7e800",
         962 => x"33676700",
         963 => x"13530501",
         964 => x"b3de6702",
         965 => x"13180501",
         966 => x"13580801",
         967 => x"93560701",
         968 => x"3316b600",
         969 => x"b3f76702",
         970 => x"330ed803",
         971 => x"93970701",
         972 => x"b3e6f600",
         973 => x"93870e00",
         974 => x"63fec601",
         975 => x"b306d500",
         976 => x"9387feff",
         977 => x"63e8a600",
         978 => x"63f6c601",
         979 => x"9387eeff",
         980 => x"b386a600",
         981 => x"b386c641",
         982 => x"33de6602",
         983 => x"13170701",
         984 => x"13570701",
         985 => x"b3f66602",
         986 => x"3308c803",
         987 => x"93960601",
         988 => x"3367d700",
         989 => x"93060e00",
         990 => x"637e0701",
         991 => x"3307e500",
         992 => x"9306feff",
         993 => x"6368a700",
         994 => x"63760701",
         995 => x"9306eeff",
         996 => x"3307a700",
         997 => x"93970701",
         998 => x"33e5d700",
         999 => x"13130601",
        1000 => x"93960601",
        1001 => x"93d60601",
        1002 => x"13530301",
        1003 => x"13560601",
        1004 => x"33070741",
        1005 => x"13580501",
        1006 => x"338e6602",
        1007 => x"33036802",
        1008 => x"93570e01",
        1009 => x"b386c602",
        1010 => x"b3866600",
        1011 => x"b387d700",
        1012 => x"3308c802",
        1013 => x"63f66700",
        1014 => x"b7060100",
        1015 => x"3308d800",
        1016 => x"93d60701",
        1017 => x"b3860601",
        1018 => x"6362d702",
        1019 => x"e31cd7ce",
        1020 => x"131e0e01",
        1021 => x"93970701",
        1022 => x"135e0e01",
        1023 => x"b398b800",
        1024 => x"b387c701",
        1025 => x"93050000",
        1026 => x"e3f0f8ce",
        1027 => x"1305f5ff",
        1028 => x"6ff05fcd",
        1029 => x"93050000",
        1030 => x"13050000",
        1031 => x"67800000",
        1032 => x"13080600",
        1033 => x"93070500",
        1034 => x"13870500",
        1035 => x"63960620",
        1036 => x"b7480000",
        1037 => x"93880896",
        1038 => x"63fcc50c",
        1039 => x"b7060100",
        1040 => x"637ed60a",
        1041 => x"93360610",
        1042 => x"93b61600",
        1043 => x"93963600",
        1044 => x"3353d600",
        1045 => x"b3886800",
        1046 => x"83c80800",
        1047 => x"13030002",
        1048 => x"b386d800",
        1049 => x"b308d340",
        1050 => x"630cd300",
        1051 => x"33971501",
        1052 => x"b356d500",
        1053 => x"33181601",
        1054 => x"33e7e600",
        1055 => x"b3171501",
        1056 => x"13560801",
        1057 => x"b356c702",
        1058 => x"13150801",
        1059 => x"13550501",
        1060 => x"3377c702",
        1061 => x"b386a602",
        1062 => x"93150701",
        1063 => x"13d70701",
        1064 => x"3367b700",
        1065 => x"637ad700",
        1066 => x"3307e800",
        1067 => x"63660701",
        1068 => x"6374d700",
        1069 => x"33070701",
        1070 => x"3307d740",
        1071 => x"b356c702",
        1072 => x"3377c702",
        1073 => x"b386a602",
        1074 => x"93970701",
        1075 => x"13170701",
        1076 => x"93d70701",
        1077 => x"b3e7e700",
        1078 => x"63fad700",
        1079 => x"b307f800",
        1080 => x"63e60701",
        1081 => x"63f4d700",
        1082 => x"b3870701",
        1083 => x"b387d740",
        1084 => x"33d51701",
        1085 => x"93050000",
        1086 => x"67800000",
        1087 => x"37030001",
        1088 => x"93068001",
        1089 => x"e37666f4",
        1090 => x"93060001",
        1091 => x"6ff05ff4",
        1092 => x"93060000",
        1093 => x"630c0600",
        1094 => x"37070100",
        1095 => x"637ee606",
        1096 => x"93360610",
        1097 => x"93b61600",
        1098 => x"93963600",
        1099 => x"3357d600",
        1100 => x"b388e800",
        1101 => x"03c70800",
        1102 => x"3307d700",
        1103 => x"93060002",
        1104 => x"b388e640",
        1105 => x"6394e606",
        1106 => x"3387c540",
        1107 => x"93550801",
        1108 => x"3356b702",
        1109 => x"13150801",
        1110 => x"13550501",
        1111 => x"93d60701",
        1112 => x"3377b702",
        1113 => x"3306a602",
        1114 => x"13170701",
        1115 => x"33e7e600",
        1116 => x"637ac700",
        1117 => x"3307e800",
        1118 => x"63660701",
        1119 => x"6374c700",
        1120 => x"33070701",
        1121 => x"3307c740",
        1122 => x"b356b702",
        1123 => x"3377b702",
        1124 => x"b386a602",
        1125 => x"6ff05ff3",
        1126 => x"37070001",
        1127 => x"93068001",
        1128 => x"e376e6f8",
        1129 => x"93060001",
        1130 => x"6ff05ff8",
        1131 => x"33181601",
        1132 => x"b3d6e500",
        1133 => x"b3171501",
        1134 => x"b3951501",
        1135 => x"3357e500",
        1136 => x"13550801",
        1137 => x"3367b700",
        1138 => x"b3d5a602",
        1139 => x"13130801",
        1140 => x"13530301",
        1141 => x"b3f6a602",
        1142 => x"b3856502",
        1143 => x"13960601",
        1144 => x"93560701",
        1145 => x"b3e6c600",
        1146 => x"63fab600",
        1147 => x"b306d800",
        1148 => x"63e60601",
        1149 => x"63f4b600",
        1150 => x"b3860601",
        1151 => x"b386b640",
        1152 => x"33d6a602",
        1153 => x"13170701",
        1154 => x"13570701",
        1155 => x"b3f6a602",
        1156 => x"33066602",
        1157 => x"93960601",
        1158 => x"3367d700",
        1159 => x"637ac700",
        1160 => x"3307e800",
        1161 => x"63660701",
        1162 => x"6374c700",
        1163 => x"33070701",
        1164 => x"3307c740",
        1165 => x"6ff09ff1",
        1166 => x"63e2d51c",
        1167 => x"37080100",
        1168 => x"63fe0605",
        1169 => x"13b80610",
        1170 => x"13381800",
        1171 => x"13183800",
        1172 => x"b7480000",
        1173 => x"33d30601",
        1174 => x"93880896",
        1175 => x"b3886800",
        1176 => x"83c80800",
        1177 => x"13030002",
        1178 => x"b3880801",
        1179 => x"33081341",
        1180 => x"63101305",
        1181 => x"63e4b600",
        1182 => x"636cc500",
        1183 => x"3306c540",
        1184 => x"b386d540",
        1185 => x"3337c500",
        1186 => x"93070600",
        1187 => x"3387e640",
        1188 => x"13850700",
        1189 => x"93050700",
        1190 => x"67800000",
        1191 => x"b7080001",
        1192 => x"13088001",
        1193 => x"e3f616fb",
        1194 => x"13080001",
        1195 => x"6ff05ffa",
        1196 => x"b3571601",
        1197 => x"b3960601",
        1198 => x"b3e6d700",
        1199 => x"33d71501",
        1200 => x"13d30601",
        1201 => x"335f6702",
        1202 => x"139e0601",
        1203 => x"135e0e01",
        1204 => x"b3970501",
        1205 => x"b3551501",
        1206 => x"b3e5f500",
        1207 => x"93d70501",
        1208 => x"33160601",
        1209 => x"33150501",
        1210 => x"33776702",
        1211 => x"b30eee03",
        1212 => x"13170701",
        1213 => x"b3e7e700",
        1214 => x"13070f00",
        1215 => x"63fed701",
        1216 => x"b387f600",
        1217 => x"1307ffff",
        1218 => x"63e8d700",
        1219 => x"63f6d701",
        1220 => x"1307efff",
        1221 => x"b387d700",
        1222 => x"b387d741",
        1223 => x"b3de6702",
        1224 => x"93950501",
        1225 => x"93d50501",
        1226 => x"b3f76702",
        1227 => x"13830e00",
        1228 => x"330ede03",
        1229 => x"93970701",
        1230 => x"b3e5f500",
        1231 => x"63fec501",
        1232 => x"b385b600",
        1233 => x"1383feff",
        1234 => x"63e8d500",
        1235 => x"63f6c501",
        1236 => x"1383eeff",
        1237 => x"b385d500",
        1238 => x"93170701",
        1239 => x"b3e76700",
        1240 => x"b385c541",
        1241 => x"13130301",
        1242 => x"131e0601",
        1243 => x"13570601",
        1244 => x"13530301",
        1245 => x"93d70701",
        1246 => x"135e0e01",
        1247 => x"b30ec303",
        1248 => x"338ec703",
        1249 => x"3303e302",
        1250 => x"b387e702",
        1251 => x"3303c301",
        1252 => x"13d70e01",
        1253 => x"33076700",
        1254 => x"6376c701",
        1255 => x"37030100",
        1256 => x"b3876700",
        1257 => x"13530701",
        1258 => x"939e0e01",
        1259 => x"13170701",
        1260 => x"93de0e01",
        1261 => x"b307f300",
        1262 => x"3307d701",
        1263 => x"63e6f500",
        1264 => x"639ef500",
        1265 => x"637ce500",
        1266 => x"3306c740",
        1267 => x"3333c700",
        1268 => x"b306d300",
        1269 => x"13070600",
        1270 => x"b387d740",
        1271 => x"3307e540",
        1272 => x"3335e500",
        1273 => x"b385f540",
        1274 => x"b385a540",
        1275 => x"b3981501",
        1276 => x"33570701",
        1277 => x"33e5e800",
        1278 => x"b3d50501",
        1279 => x"67800000",
        1280 => x"13030500",
        1281 => x"630a0600",
        1282 => x"2300b300",
        1283 => x"1306f6ff",
        1284 => x"13031300",
        1285 => x"e31a06fe",
        1286 => x"67800000",
        1287 => x"13030500",
        1288 => x"630e0600",
        1289 => x"83830500",
        1290 => x"23007300",
        1291 => x"1306f6ff",
        1292 => x"13031300",
        1293 => x"93851500",
        1294 => x"e31606fe",
        1295 => x"67800000",
        1296 => x"630c0602",
        1297 => x"13030500",
        1298 => x"93061000",
        1299 => x"636ab500",
        1300 => x"9306f0ff",
        1301 => x"1307f6ff",
        1302 => x"3303e300",
        1303 => x"b385e500",
        1304 => x"83830500",
        1305 => x"23007300",
        1306 => x"1306f6ff",
        1307 => x"3303d300",
        1308 => x"b385d500",
        1309 => x"e31606fe",
        1310 => x"67800000",
        1311 => x"370700f0",
        1312 => x"13070710",
        1313 => x"83274700",
        1314 => x"93f78700",
        1315 => x"e38c07fe",
        1316 => x"03258700",
        1317 => x"1375f50f",
        1318 => x"67800000",
        1319 => x"f32710fc",
        1320 => x"63960700",
        1321 => x"b7f7fa02",
        1322 => x"93870708",
        1323 => x"63060500",
        1324 => x"33d5a702",
        1325 => x"1305f5ff",
        1326 => x"b70700f0",
        1327 => x"23a6a710",
        1328 => x"23a0b710",
        1329 => x"23a20710",
        1330 => x"67800000",
        1331 => x"370700f0",
        1332 => x"1375f50f",
        1333 => x"13070710",
        1334 => x"2324a700",
        1335 => x"83274700",
        1336 => x"93f70701",
        1337 => x"e38c07fe",
        1338 => x"67800000",
        1339 => x"630e0502",
        1340 => x"130101ff",
        1341 => x"23248100",
        1342 => x"23261100",
        1343 => x"13040500",
        1344 => x"03450500",
        1345 => x"630a0500",
        1346 => x"13041400",
        1347 => x"eff01ffc",
        1348 => x"03450400",
        1349 => x"e31a05fe",
        1350 => x"8320c100",
        1351 => x"03248100",
        1352 => x"13010101",
        1353 => x"67800000",
        1354 => x"67800000",
        1355 => x"130101f9",
        1356 => x"23229106",
        1357 => x"23202107",
        1358 => x"23261106",
        1359 => x"23248106",
        1360 => x"232e3105",
        1361 => x"232c4105",
        1362 => x"232a5105",
        1363 => x"23286105",
        1364 => x"23267105",
        1365 => x"23248105",
        1366 => x"23229105",
        1367 => x"13090500",
        1368 => x"93840500",
        1369 => x"f32a00fc",
        1370 => x"b7070008",
        1371 => x"232c0100",
        1372 => x"232e0100",
        1373 => x"23200102",
        1374 => x"23220102",
        1375 => x"23240102",
        1376 => x"23260102",
        1377 => x"23280102",
        1378 => x"232a0102",
        1379 => x"232c0102",
        1380 => x"232e0102",
        1381 => x"b3fafa00",
        1382 => x"732410fc",
        1383 => x"63160400",
        1384 => x"37f4fa02",
        1385 => x"13040408",
        1386 => x"97f2ffff",
        1387 => x"938282d5",
        1388 => x"73905230",
        1389 => x"37c50100",
        1390 => x"13050520",
        1391 => x"93059000",
        1392 => x"eff0dfed",
        1393 => x"b717b7d1",
        1394 => x"93879775",
        1395 => x"b337f402",
        1396 => x"93561400",
        1397 => x"37353e05",
        1398 => x"370600f0",
        1399 => x"13576400",
        1400 => x"130535d6",
        1401 => x"9386f6ff",
        1402 => x"2326d660",
        1403 => x"b725d96f",
        1404 => x"93060600",
        1405 => x"3337a702",
        1406 => x"93d7d700",
        1407 => x"13051001",
        1408 => x"2320a660",
        1409 => x"938555d8",
        1410 => x"9387f7ff",
        1411 => x"23a8f670",
        1412 => x"37260000",
        1413 => x"1306f670",
        1414 => x"23a6c670",
        1415 => x"b337b402",
        1416 => x"13576700",
        1417 => x"1307f7ff",
        1418 => x"23a0a670",
        1419 => x"93058070",
        1420 => x"13170701",
        1421 => x"23a0b640",
        1422 => x"13678700",
        1423 => x"23a0e620",
        1424 => x"1307a007",
        1425 => x"93d73701",
        1426 => x"9387f7ff",
        1427 => x"93970701",
        1428 => x"93e7c700",
        1429 => x"23a0f630",
        1430 => x"23ace600",
        1431 => x"f3224030",
        1432 => x"93e20208",
        1433 => x"73904230",
        1434 => x"f3224030",
        1435 => x"93e28200",
        1436 => x"73904230",
        1437 => x"b7220000",
        1438 => x"93828280",
        1439 => x"73900230",
        1440 => x"b7490000",
        1441 => x"138509a8",
        1442 => x"eff05fe6",
        1443 => x"1304f9ff",
        1444 => x"63522003",
        1445 => x"1309f0ff",
        1446 => x"03a50400",
        1447 => x"1304f4ff",
        1448 => x"93844400",
        1449 => x"eff09fe4",
        1450 => x"138509a8",
        1451 => x"eff01fe4",
        1452 => x"e31424ff",
        1453 => x"37450000",
        1454 => x"130545a8",
        1455 => x"eff01fe3",
        1456 => x"63960a22",
        1457 => x"b7040010",
        1458 => x"b7998888",
        1459 => x"37f4eeee",
        1460 => x"9384f4ff",
        1461 => x"93899988",
        1462 => x"1304f4ee",
        1463 => x"374a0000",
        1464 => x"b71b0000",
        1465 => x"37f9eeee",
        1466 => x"938b0b2c",
        1467 => x"1309e9ee",
        1468 => x"6f00c000",
        1469 => x"938bfbff",
        1470 => x"63860b1a",
        1471 => x"93050000",
        1472 => x"13058100",
        1473 => x"ef00d030",
        1474 => x"e31605fe",
        1475 => x"032c8100",
        1476 => x"8325c100",
        1477 => x"37160000",
        1478 => x"9357cc01",
        1479 => x"13974500",
        1480 => x"b367f700",
        1481 => x"33f79700",
        1482 => x"b3779c00",
        1483 => x"13d58501",
        1484 => x"b387e700",
        1485 => x"13d7f541",
        1486 => x"b387a700",
        1487 => x"1375d700",
        1488 => x"b387a700",
        1489 => x"33b83703",
        1490 => x"137727ff",
        1491 => x"130606e1",
        1492 => x"93060000",
        1493 => x"13050c00",
        1494 => x"938bfbff",
        1495 => x"13583800",
        1496 => x"93184800",
        1497 => x"33880841",
        1498 => x"b3870741",
        1499 => x"b387e700",
        1500 => x"13d7f741",
        1501 => x"b307fc40",
        1502 => x"3338fc00",
        1503 => x"3387e540",
        1504 => x"33070741",
        1505 => x"b3882703",
        1506 => x"33078702",
        1507 => x"33b88702",
        1508 => x"33071701",
        1509 => x"b3878702",
        1510 => x"33070701",
        1511 => x"1358f741",
        1512 => x"13783800",
        1513 => x"b307f800",
        1514 => x"33b80701",
        1515 => x"3308e800",
        1516 => x"1317e801",
        1517 => x"93d72700",
        1518 => x"b367f700",
        1519 => x"93582840",
        1520 => x"13d7c701",
        1521 => x"13934800",
        1522 => x"3367e300",
        1523 => x"33739700",
        1524 => x"33f79700",
        1525 => x"1358f841",
        1526 => x"33076700",
        1527 => x"13d38801",
        1528 => x"33076700",
        1529 => x"1373d800",
        1530 => x"33076700",
        1531 => x"33333703",
        1532 => x"137828ff",
        1533 => x"139b4700",
        1534 => x"330bfb40",
        1535 => x"131b2b00",
        1536 => x"330b6c41",
        1537 => x"13533300",
        1538 => x"131e4300",
        1539 => x"33036e40",
        1540 => x"33076740",
        1541 => x"33070701",
        1542 => x"1358f741",
        1543 => x"3387e740",
        1544 => x"33880841",
        1545 => x"b3b8e700",
        1546 => x"33081841",
        1547 => x"33032703",
        1548 => x"33088802",
        1549 => x"b3388702",
        1550 => x"33086800",
        1551 => x"33078702",
        1552 => x"33081801",
        1553 => x"9358f841",
        1554 => x"93f83800",
        1555 => x"3387e800",
        1556 => x"b3381701",
        1557 => x"b3880801",
        1558 => x"9398e801",
        1559 => x"13572700",
        1560 => x"33e7e800",
        1561 => x"13184700",
        1562 => x"3307e840",
        1563 => x"13172700",
        1564 => x"b38ce740",
        1565 => x"efe0dff0",
        1566 => x"83260101",
        1567 => x"13070500",
        1568 => x"13080b00",
        1569 => x"93870c00",
        1570 => x"13060c00",
        1571 => x"9305caae",
        1572 => x"13058101",
        1573 => x"ef008047",
        1574 => x"13058101",
        1575 => x"eff01fc5",
        1576 => x"e39e0be4",
        1577 => x"63940a00",
        1578 => x"73001000",
        1579 => x"b70700f0",
        1580 => x"9306f00f",
        1581 => x"23a4d740",
        1582 => x"83a60720",
        1583 => x"13060009",
        1584 => x"371700f0",
        1585 => x"93e60630",
        1586 => x"23a0d720",
        1587 => x"23a4c720",
        1588 => x"83a60730",
        1589 => x"93e60630",
        1590 => x"23a0d730",
        1591 => x"23a4c730",
        1592 => x"93071000",
        1593 => x"2320f790",
        1594 => x"6ff09fdf",
        1595 => x"37450000",
        1596 => x"130545ab",
        1597 => x"eff09fbf",
        1598 => x"6ff0dfdc",
        1599 => x"130101ff",
        1600 => x"23248100",
        1601 => x"23261100",
        1602 => x"93070000",
        1603 => x"13040500",
        1604 => x"63880700",
        1605 => x"93050000",
        1606 => x"97000000",
        1607 => x"e7000000",
        1608 => x"83a74187",
        1609 => x"63840700",
        1610 => x"e7800700",
        1611 => x"13050400",
        1612 => x"ef101047",
        1613 => x"13050000",
        1614 => x"67800000",
        1615 => x"130101ff",
        1616 => x"23248100",
        1617 => x"23261100",
        1618 => x"13040500",
        1619 => x"2316b500",
        1620 => x"2317c500",
        1621 => x"23200500",
        1622 => x"23220500",
        1623 => x"23240500",
        1624 => x"23220506",
        1625 => x"23280500",
        1626 => x"232a0500",
        1627 => x"232c0500",
        1628 => x"13068000",
        1629 => x"93050000",
        1630 => x"1305c505",
        1631 => x"eff05fa8",
        1632 => x"b7270000",
        1633 => x"938707d8",
        1634 => x"2322f402",
        1635 => x"b7270000",
        1636 => x"938787dd",
        1637 => x"2324f402",
        1638 => x"b7270000",
        1639 => x"9387c7e5",
        1640 => x"2326f402",
        1641 => x"b7270000",
        1642 => x"938747eb",
        1643 => x"8320c100",
        1644 => x"23208402",
        1645 => x"2328f402",
        1646 => x"03248100",
        1647 => x"13010101",
        1648 => x"67800000",
        1649 => x"b7350000",
        1650 => x"37050020",
        1651 => x"13868181",
        1652 => x"93854532",
        1653 => x"13054502",
        1654 => x"6f00c021",
        1655 => x"83254500",
        1656 => x"130101ff",
        1657 => x"b7070020",
        1658 => x"23248100",
        1659 => x"23261100",
        1660 => x"93878708",
        1661 => x"13040500",
        1662 => x"6384f500",
        1663 => x"ef109012",
        1664 => x"83258400",
        1665 => x"9387018f",
        1666 => x"6386f500",
        1667 => x"13050400",
        1668 => x"ef105011",
        1669 => x"8325c400",
        1670 => x"93878195",
        1671 => x"638cf500",
        1672 => x"13050400",
        1673 => x"03248100",
        1674 => x"8320c100",
        1675 => x"13010101",
        1676 => x"6f10500f",
        1677 => x"8320c100",
        1678 => x"03248100",
        1679 => x"13010101",
        1680 => x"67800000",
        1681 => x"b7270000",
        1682 => x"37050020",
        1683 => x"130101ff",
        1684 => x"9387479c",
        1685 => x"13060000",
        1686 => x"93054000",
        1687 => x"13058508",
        1688 => x"23261100",
        1689 => x"23aaf186",
        1690 => x"eff05fed",
        1691 => x"13061000",
        1692 => x"93059000",
        1693 => x"1385018f",
        1694 => x"eff05fec",
        1695 => x"8320c100",
        1696 => x"13062000",
        1697 => x"93052001",
        1698 => x"13858195",
        1699 => x"13010101",
        1700 => x"6ff0dfea",
        1701 => x"13050000",
        1702 => x"67800000",
        1703 => x"83a74187",
        1704 => x"130101ff",
        1705 => x"23202101",
        1706 => x"23261100",
        1707 => x"23248100",
        1708 => x"23229100",
        1709 => x"13090500",
        1710 => x"63940700",
        1711 => x"eff09ff8",
        1712 => x"93848181",
        1713 => x"03a48400",
        1714 => x"83a74400",
        1715 => x"9387f7ff",
        1716 => x"63d80702",
        1717 => x"03a40400",
        1718 => x"6310040c",
        1719 => x"9305c01a",
        1720 => x"13050900",
        1721 => x"ef00900b",
        1722 => x"13040500",
        1723 => x"63140508",
        1724 => x"23a00400",
        1725 => x"9307c000",
        1726 => x"2320f900",
        1727 => x"6f004005",
        1728 => x"0317c400",
        1729 => x"63140706",
        1730 => x"b707ffff",
        1731 => x"93871700",
        1732 => x"23220406",
        1733 => x"23200400",
        1734 => x"23220400",
        1735 => x"23240400",
        1736 => x"2326f400",
        1737 => x"23280400",
        1738 => x"232a0400",
        1739 => x"232c0400",
        1740 => x"13068000",
        1741 => x"93050000",
        1742 => x"1305c405",
        1743 => x"eff05f8c",
        1744 => x"232a0402",
        1745 => x"232c0402",
        1746 => x"23240404",
        1747 => x"23260404",
        1748 => x"8320c100",
        1749 => x"13050400",
        1750 => x"03248100",
        1751 => x"83244100",
        1752 => x"03290100",
        1753 => x"13010101",
        1754 => x"67800000",
        1755 => x"13048406",
        1756 => x"6ff0dff5",
        1757 => x"93074000",
        1758 => x"23200500",
        1759 => x"2322f500",
        1760 => x"1305c500",
        1761 => x"2324a400",
        1762 => x"1306001a",
        1763 => x"93050000",
        1764 => x"eff01f87",
        1765 => x"23a08400",
        1766 => x"93040400",
        1767 => x"6ff09ff2",
        1768 => x"83270502",
        1769 => x"639e0700",
        1770 => x"b7270000",
        1771 => x"9387c79d",
        1772 => x"2320f502",
        1773 => x"83a74187",
        1774 => x"63940700",
        1775 => x"6ff09fe8",
        1776 => x"67800000",
        1777 => x"67800000",
        1778 => x"67800000",
        1779 => x"b7250000",
        1780 => x"13868181",
        1781 => x"93854593",
        1782 => x"13050000",
        1783 => x"6f008001",
        1784 => x"b7250000",
        1785 => x"13868181",
        1786 => x"938545a9",
        1787 => x"13050000",
        1788 => x"6f004000",
        1789 => x"130101fd",
        1790 => x"23248102",
        1791 => x"23202103",
        1792 => x"232e3101",
        1793 => x"232c4101",
        1794 => x"23286101",
        1795 => x"23267101",
        1796 => x"23261102",
        1797 => x"23229102",
        1798 => x"232a5101",
        1799 => x"93090500",
        1800 => x"138a0500",
        1801 => x"13040600",
        1802 => x"13090000",
        1803 => x"130b1000",
        1804 => x"930bf0ff",
        1805 => x"83248400",
        1806 => x"832a4400",
        1807 => x"938afaff",
        1808 => x"63de0a02",
        1809 => x"03240400",
        1810 => x"e31604fe",
        1811 => x"8320c102",
        1812 => x"03248102",
        1813 => x"83244102",
        1814 => x"8329c101",
        1815 => x"032a8101",
        1816 => x"832a4101",
        1817 => x"032b0101",
        1818 => x"832bc100",
        1819 => x"13050900",
        1820 => x"03290102",
        1821 => x"13010103",
        1822 => x"67800000",
        1823 => x"83d7c400",
        1824 => x"637efb00",
        1825 => x"8397e400",
        1826 => x"638a7701",
        1827 => x"93850400",
        1828 => x"13850900",
        1829 => x"e7000a00",
        1830 => x"3369a900",
        1831 => x"93848406",
        1832 => x"6ff0dff9",
        1833 => x"130101f6",
        1834 => x"232af108",
        1835 => x"b7070080",
        1836 => x"9387f7ff",
        1837 => x"232ef100",
        1838 => x"2328f100",
        1839 => x"b707ffff",
        1840 => x"2326d108",
        1841 => x"2324b100",
        1842 => x"232cb100",
        1843 => x"93878720",
        1844 => x"9306c108",
        1845 => x"93058100",
        1846 => x"232e1106",
        1847 => x"232af100",
        1848 => x"2328e108",
        1849 => x"232c0109",
        1850 => x"232e1109",
        1851 => x"23260106",
        1852 => x"2322d100",
        1853 => x"ef00103a",
        1854 => x"83278100",
        1855 => x"23800700",
        1856 => x"8320c107",
        1857 => x"1301010a",
        1858 => x"67800000",
        1859 => x"130101f6",
        1860 => x"232af108",
        1861 => x"b7070080",
        1862 => x"9387f7ff",
        1863 => x"232ef100",
        1864 => x"2328f100",
        1865 => x"b707ffff",
        1866 => x"93878720",
        1867 => x"232af100",
        1868 => x"2324a100",
        1869 => x"232ca100",
        1870 => x"03a50187",
        1871 => x"2324c108",
        1872 => x"2326d108",
        1873 => x"13860500",
        1874 => x"93068108",
        1875 => x"93058100",
        1876 => x"232e1106",
        1877 => x"2328e108",
        1878 => x"232c0109",
        1879 => x"232e1109",
        1880 => x"23260106",
        1881 => x"2322d100",
        1882 => x"ef00d032",
        1883 => x"83278100",
        1884 => x"23800700",
        1885 => x"8320c107",
        1886 => x"1301010a",
        1887 => x"67800000",
        1888 => x"130101ff",
        1889 => x"23248100",
        1890 => x"13840500",
        1891 => x"8395e500",
        1892 => x"23261100",
        1893 => x"ef008033",
        1894 => x"63400502",
        1895 => x"83274405",
        1896 => x"b387a700",
        1897 => x"232af404",
        1898 => x"8320c100",
        1899 => x"03248100",
        1900 => x"13010101",
        1901 => x"67800000",
        1902 => x"8357c400",
        1903 => x"37f7ffff",
        1904 => x"1307f7ff",
        1905 => x"b3f7e700",
        1906 => x"2316f400",
        1907 => x"6ff0dffd",
        1908 => x"13050000",
        1909 => x"67800000",
        1910 => x"83d7c500",
        1911 => x"130101fe",
        1912 => x"232c8100",
        1913 => x"232a9100",
        1914 => x"23282101",
        1915 => x"23263101",
        1916 => x"232e1100",
        1917 => x"93f70710",
        1918 => x"93040500",
        1919 => x"13840500",
        1920 => x"13090600",
        1921 => x"93890600",
        1922 => x"638a0700",
        1923 => x"8395e500",
        1924 => x"93062000",
        1925 => x"13060000",
        1926 => x"ef004026",
        1927 => x"8357c400",
        1928 => x"37f7ffff",
        1929 => x"1307f7ff",
        1930 => x"b3f7e700",
        1931 => x"8315e400",
        1932 => x"2316f400",
        1933 => x"03248101",
        1934 => x"8320c101",
        1935 => x"93860900",
        1936 => x"13060900",
        1937 => x"8329c100",
        1938 => x"03290101",
        1939 => x"13850400",
        1940 => x"83244101",
        1941 => x"13010102",
        1942 => x"6f00402c",
        1943 => x"130101ff",
        1944 => x"23248100",
        1945 => x"13840500",
        1946 => x"8395e500",
        1947 => x"23261100",
        1948 => x"ef00c020",
        1949 => x"1307f0ff",
        1950 => x"8317c400",
        1951 => x"6312e502",
        1952 => x"37f7ffff",
        1953 => x"1307f7ff",
        1954 => x"b3f7e700",
        1955 => x"2316f400",
        1956 => x"8320c100",
        1957 => x"03248100",
        1958 => x"13010101",
        1959 => x"67800000",
        1960 => x"37170000",
        1961 => x"b3e7e700",
        1962 => x"2316f400",
        1963 => x"232aa404",
        1964 => x"6ff01ffe",
        1965 => x"8395e500",
        1966 => x"6f004000",
        1967 => x"130101ff",
        1968 => x"23248100",
        1969 => x"23229100",
        1970 => x"13040500",
        1971 => x"13850500",
        1972 => x"23261100",
        1973 => x"23ac0186",
        1974 => x"ef108068",
        1975 => x"9307f0ff",
        1976 => x"6318f500",
        1977 => x"83a78187",
        1978 => x"63840700",
        1979 => x"2320f400",
        1980 => x"8320c100",
        1981 => x"03248100",
        1982 => x"83244100",
        1983 => x"13010101",
        1984 => x"67800000",
        1985 => x"83a70187",
        1986 => x"6388a716",
        1987 => x"8327c501",
        1988 => x"130101fe",
        1989 => x"232c8100",
        1990 => x"232e1100",
        1991 => x"232a9100",
        1992 => x"23282101",
        1993 => x"23263101",
        1994 => x"13040500",
        1995 => x"63840708",
        1996 => x"83a7c700",
        1997 => x"638c0702",
        1998 => x"93040000",
        1999 => x"13090008",
        2000 => x"8327c401",
        2001 => x"83a7c700",
        2002 => x"b3879700",
        2003 => x"83a50700",
        2004 => x"63980504",
        2005 => x"93844400",
        2006 => x"e39424ff",
        2007 => x"8327c401",
        2008 => x"13050400",
        2009 => x"83a5c700",
        2010 => x"ef00802b",
        2011 => x"8327c401",
        2012 => x"83a50700",
        2013 => x"63860500",
        2014 => x"13050400",
        2015 => x"ef00402a",
        2016 => x"8327c401",
        2017 => x"83a48700",
        2018 => x"63860402",
        2019 => x"93850400",
        2020 => x"13050400",
        2021 => x"83a40400",
        2022 => x"ef008028",
        2023 => x"6ff0dffe",
        2024 => x"83a90500",
        2025 => x"13050400",
        2026 => x"ef008027",
        2027 => x"93850900",
        2028 => x"6ff01ffa",
        2029 => x"83254401",
        2030 => x"63860500",
        2031 => x"13050400",
        2032 => x"ef000026",
        2033 => x"8325c401",
        2034 => x"63860500",
        2035 => x"13050400",
        2036 => x"ef000025",
        2037 => x"83250403",
        2038 => x"63860500",
        2039 => x"13050400",
        2040 => x"ef000024",
        2041 => x"83254403",
        2042 => x"63860500",
        2043 => x"13050400",
        2044 => x"ef000023",
        2045 => x"83258403",
        2046 => x"63860500",
        2047 => x"13050400",
        2048 => x"ef000022",
        2049 => x"83258404",
        2050 => x"63860500",
        2051 => x"13050400",
        2052 => x"ef000021",
        2053 => x"83254404",
        2054 => x"63860500",
        2055 => x"13050400",
        2056 => x"ef000020",
        2057 => x"8325c402",
        2058 => x"63860500",
        2059 => x"13050400",
        2060 => x"ef00001f",
        2061 => x"83270402",
        2062 => x"63820702",
        2063 => x"13050400",
        2064 => x"03248101",
        2065 => x"8320c101",
        2066 => x"83244101",
        2067 => x"03290101",
        2068 => x"8329c100",
        2069 => x"13010102",
        2070 => x"67800700",
        2071 => x"8320c101",
        2072 => x"03248101",
        2073 => x"83244101",
        2074 => x"03290101",
        2075 => x"8329c100",
        2076 => x"13010102",
        2077 => x"67800000",
        2078 => x"67800000",
        2079 => x"130101ff",
        2080 => x"23248100",
        2081 => x"23229100",
        2082 => x"13040500",
        2083 => x"13850500",
        2084 => x"93050600",
        2085 => x"13860600",
        2086 => x"23261100",
        2087 => x"23ac0186",
        2088 => x"ef10405a",
        2089 => x"9307f0ff",
        2090 => x"6318f500",
        2091 => x"83a78187",
        2092 => x"63840700",
        2093 => x"2320f400",
        2094 => x"8320c100",
        2095 => x"03248100",
        2096 => x"83244100",
        2097 => x"13010101",
        2098 => x"67800000",
        2099 => x"130101ff",
        2100 => x"23248100",
        2101 => x"23229100",
        2102 => x"13040500",
        2103 => x"13850500",
        2104 => x"93050600",
        2105 => x"13860600",
        2106 => x"23261100",
        2107 => x"23ac0186",
        2108 => x"ef104059",
        2109 => x"9307f0ff",
        2110 => x"6318f500",
        2111 => x"83a78187",
        2112 => x"63840700",
        2113 => x"2320f400",
        2114 => x"8320c100",
        2115 => x"03248100",
        2116 => x"83244100",
        2117 => x"13010101",
        2118 => x"67800000",
        2119 => x"130101ff",
        2120 => x"23248100",
        2121 => x"23229100",
        2122 => x"13040500",
        2123 => x"13850500",
        2124 => x"93050600",
        2125 => x"13860600",
        2126 => x"23261100",
        2127 => x"23ac0186",
        2128 => x"ef10c05e",
        2129 => x"9307f0ff",
        2130 => x"6318f500",
        2131 => x"83a78187",
        2132 => x"63840700",
        2133 => x"2320f400",
        2134 => x"8320c100",
        2135 => x"03248100",
        2136 => x"83244100",
        2137 => x"13010101",
        2138 => x"67800000",
        2139 => x"03a50187",
        2140 => x"67800000",
        2141 => x"130101ff",
        2142 => x"23248100",
        2143 => x"23229100",
        2144 => x"37440000",
        2145 => x"b7440000",
        2146 => x"9387c4c4",
        2147 => x"1304c4c4",
        2148 => x"3304f440",
        2149 => x"23202101",
        2150 => x"23261100",
        2151 => x"13542440",
        2152 => x"9384c4c4",
        2153 => x"13090000",
        2154 => x"63108904",
        2155 => x"b7440000",
        2156 => x"37440000",
        2157 => x"9387c4c4",
        2158 => x"1304c4c4",
        2159 => x"3304f440",
        2160 => x"13542440",
        2161 => x"9384c4c4",
        2162 => x"13090000",
        2163 => x"63188902",
        2164 => x"8320c100",
        2165 => x"03248100",
        2166 => x"83244100",
        2167 => x"03290100",
        2168 => x"13010101",
        2169 => x"67800000",
        2170 => x"83a70400",
        2171 => x"13091900",
        2172 => x"93844400",
        2173 => x"e7800700",
        2174 => x"6ff01ffb",
        2175 => x"83a70400",
        2176 => x"13091900",
        2177 => x"93844400",
        2178 => x"e7800700",
        2179 => x"6ff01ffc",
        2180 => x"13860500",
        2181 => x"93050500",
        2182 => x"03a50187",
        2183 => x"6f10c01b",
        2184 => x"638a050e",
        2185 => x"83a7c5ff",
        2186 => x"130101fe",
        2187 => x"232c8100",
        2188 => x"232e1100",
        2189 => x"1384c5ff",
        2190 => x"63d40700",
        2191 => x"3304f400",
        2192 => x"2326a100",
        2193 => x"ef004031",
        2194 => x"83a70188",
        2195 => x"0325c100",
        2196 => x"639e0700",
        2197 => x"23220400",
        2198 => x"23a08188",
        2199 => x"03248101",
        2200 => x"8320c101",
        2201 => x"13010102",
        2202 => x"6f00402f",
        2203 => x"6374f402",
        2204 => x"03260400",
        2205 => x"b306c400",
        2206 => x"639ad700",
        2207 => x"83a60700",
        2208 => x"83a74700",
        2209 => x"b386c600",
        2210 => x"2320d400",
        2211 => x"2322f400",
        2212 => x"6ff09ffc",
        2213 => x"13870700",
        2214 => x"83a74700",
        2215 => x"63840700",
        2216 => x"e37af4fe",
        2217 => x"83260700",
        2218 => x"3306d700",
        2219 => x"63188602",
        2220 => x"03260400",
        2221 => x"b386c600",
        2222 => x"2320d700",
        2223 => x"3306d700",
        2224 => x"e39ec7f8",
        2225 => x"03a60700",
        2226 => x"83a74700",
        2227 => x"b306d600",
        2228 => x"2320d700",
        2229 => x"2322f700",
        2230 => x"6ff05ff8",
        2231 => x"6378c400",
        2232 => x"9307c000",
        2233 => x"2320f500",
        2234 => x"6ff05ff7",
        2235 => x"03260400",
        2236 => x"b306c400",
        2237 => x"639ad700",
        2238 => x"83a60700",
        2239 => x"83a74700",
        2240 => x"b386c600",
        2241 => x"2320d400",
        2242 => x"2322f400",
        2243 => x"23228700",
        2244 => x"6ff0dff4",
        2245 => x"67800000",
        2246 => x"130101ff",
        2247 => x"23202101",
        2248 => x"83a7c187",
        2249 => x"23248100",
        2250 => x"23229100",
        2251 => x"23261100",
        2252 => x"93040500",
        2253 => x"13840500",
        2254 => x"63980700",
        2255 => x"93050000",
        2256 => x"ef10400e",
        2257 => x"23aea186",
        2258 => x"93050400",
        2259 => x"13850400",
        2260 => x"ef10400d",
        2261 => x"1309f0ff",
        2262 => x"63122503",
        2263 => x"1304f0ff",
        2264 => x"8320c100",
        2265 => x"13050400",
        2266 => x"03248100",
        2267 => x"83244100",
        2268 => x"03290100",
        2269 => x"13010101",
        2270 => x"67800000",
        2271 => x"13043500",
        2272 => x"1374c4ff",
        2273 => x"e30e85fc",
        2274 => x"b305a440",
        2275 => x"13850400",
        2276 => x"ef104009",
        2277 => x"e31625fd",
        2278 => x"6ff05ffc",
        2279 => x"130101fe",
        2280 => x"232a9100",
        2281 => x"93843500",
        2282 => x"93f4c4ff",
        2283 => x"23282101",
        2284 => x"232e1100",
        2285 => x"232c8100",
        2286 => x"23263101",
        2287 => x"23244101",
        2288 => x"93848400",
        2289 => x"9307c000",
        2290 => x"13090500",
        2291 => x"63fef408",
        2292 => x"93840700",
        2293 => x"63ecb408",
        2294 => x"13050900",
        2295 => x"ef00c017",
        2296 => x"83a70188",
        2297 => x"13840700",
        2298 => x"6316040a",
        2299 => x"93850400",
        2300 => x"13050900",
        2301 => x"eff05ff2",
        2302 => x"9307f0ff",
        2303 => x"13040500",
        2304 => x"6318f514",
        2305 => x"03a40188",
        2306 => x"93070400",
        2307 => x"63980710",
        2308 => x"63060412",
        2309 => x"032a0400",
        2310 => x"93050000",
        2311 => x"13050900",
        2312 => x"330a4401",
        2313 => x"ef100000",
        2314 => x"631aaa10",
        2315 => x"83270400",
        2316 => x"13050900",
        2317 => x"b384f440",
        2318 => x"93850400",
        2319 => x"eff0dfed",
        2320 => x"9307f0ff",
        2321 => x"630cf50e",
        2322 => x"83270400",
        2323 => x"b3879700",
        2324 => x"2320f400",
        2325 => x"83a70188",
        2326 => x"03a74700",
        2327 => x"6316070c",
        2328 => x"23a00188",
        2329 => x"6f000006",
        2330 => x"e3d604f6",
        2331 => x"2320f900",
        2332 => x"13050000",
        2333 => x"8320c101",
        2334 => x"03248101",
        2335 => x"83244101",
        2336 => x"03290101",
        2337 => x"8329c100",
        2338 => x"032a8100",
        2339 => x"13010102",
        2340 => x"67800000",
        2341 => x"83260400",
        2342 => x"b3869640",
        2343 => x"63ca0606",
        2344 => x"1307b000",
        2345 => x"637ad704",
        2346 => x"23209400",
        2347 => x"33079400",
        2348 => x"63908704",
        2349 => x"23a0e188",
        2350 => x"83274400",
        2351 => x"2320d700",
        2352 => x"2322f700",
        2353 => x"13050900",
        2354 => x"ef004009",
        2355 => x"1305b400",
        2356 => x"93074400",
        2357 => x"137585ff",
        2358 => x"3307f540",
        2359 => x"e30cf5f8",
        2360 => x"3304e400",
        2361 => x"b387a740",
        2362 => x"2320f400",
        2363 => x"6ff09ff8",
        2364 => x"23a2e700",
        2365 => x"6ff05ffc",
        2366 => x"03274400",
        2367 => x"63968700",
        2368 => x"23a0e188",
        2369 => x"6ff01ffc",
        2370 => x"23a2e700",
        2371 => x"6ff09ffb",
        2372 => x"93070400",
        2373 => x"03244400",
        2374 => x"6ff01fed",
        2375 => x"13840700",
        2376 => x"83a74700",
        2377 => x"6ff09fee",
        2378 => x"13870700",
        2379 => x"83a74700",
        2380 => x"e39c87fe",
        2381 => x"23220700",
        2382 => x"6ff0dff8",
        2383 => x"9307c000",
        2384 => x"2320f900",
        2385 => x"13050900",
        2386 => x"ef004001",
        2387 => x"6ff05ff2",
        2388 => x"23209500",
        2389 => x"6ff01ff7",
        2390 => x"67800000",
        2391 => x"67800000",
        2392 => x"130101fe",
        2393 => x"23282101",
        2394 => x"03a98500",
        2395 => x"232c8100",
        2396 => x"23263101",
        2397 => x"23244101",
        2398 => x"232e1100",
        2399 => x"232a9100",
        2400 => x"23225101",
        2401 => x"23206101",
        2402 => x"13840500",
        2403 => x"130a0600",
        2404 => x"93890600",
        2405 => x"63ec2613",
        2406 => x"8397c500",
        2407 => x"13070900",
        2408 => x"93f60748",
        2409 => x"638c0608",
        2410 => x"83244401",
        2411 => x"13073000",
        2412 => x"83a50501",
        2413 => x"b384e402",
        2414 => x"13072000",
        2415 => x"832a0400",
        2416 => x"130b0500",
        2417 => x"b38aba40",
        2418 => x"b3c4e402",
        2419 => x"13871900",
        2420 => x"33075701",
        2421 => x"13860400",
        2422 => x"63f6e400",
        2423 => x"93040700",
        2424 => x"13060700",
        2425 => x"93f70740",
        2426 => x"6386070a",
        2427 => x"93050600",
        2428 => x"13050b00",
        2429 => x"eff09fda",
        2430 => x"13090500",
        2431 => x"630a050a",
        2432 => x"83250401",
        2433 => x"13860a00",
        2434 => x"efe05fe1",
        2435 => x"8357c400",
        2436 => x"93f7f7b7",
        2437 => x"93e70708",
        2438 => x"2316f400",
        2439 => x"23282401",
        2440 => x"232a9400",
        2441 => x"33095901",
        2442 => x"b3845441",
        2443 => x"23202401",
        2444 => x"23249400",
        2445 => x"13890900",
        2446 => x"13870900",
        2447 => x"93090700",
        2448 => x"03250400",
        2449 => x"13860900",
        2450 => x"93050a00",
        2451 => x"efe05fdf",
        2452 => x"83278400",
        2453 => x"13050000",
        2454 => x"b3872741",
        2455 => x"2324f400",
        2456 => x"83270400",
        2457 => x"b3873701",
        2458 => x"2320f400",
        2459 => x"8320c101",
        2460 => x"03248101",
        2461 => x"83244101",
        2462 => x"03290101",
        2463 => x"8329c100",
        2464 => x"032a8100",
        2465 => x"832a4100",
        2466 => x"032b0100",
        2467 => x"13010102",
        2468 => x"67800000",
        2469 => x"13050b00",
        2470 => x"ef00505d",
        2471 => x"13090500",
        2472 => x"e31e05f6",
        2473 => x"83250401",
        2474 => x"13050b00",
        2475 => x"eff05fb7",
        2476 => x"9307c000",
        2477 => x"2320fb00",
        2478 => x"8357c400",
        2479 => x"1305f0ff",
        2480 => x"93e70704",
        2481 => x"2316f400",
        2482 => x"6ff05ffa",
        2483 => x"13890600",
        2484 => x"6ff01ff7",
        2485 => x"83278600",
        2486 => x"130101fd",
        2487 => x"232e3101",
        2488 => x"23261102",
        2489 => x"23248102",
        2490 => x"23229102",
        2491 => x"23202103",
        2492 => x"232c4101",
        2493 => x"232a5101",
        2494 => x"23286101",
        2495 => x"23267101",
        2496 => x"23248101",
        2497 => x"23229101",
        2498 => x"2320a101",
        2499 => x"93090600",
        2500 => x"63800710",
        2501 => x"832a0600",
        2502 => x"130a0500",
        2503 => x"13840500",
        2504 => x"930b3000",
        2505 => x"130c2000",
        2506 => x"03ad4a00",
        2507 => x"03ab0a00",
        2508 => x"938a8a00",
        2509 => x"e30a0dfe",
        2510 => x"03298400",
        2511 => x"93040900",
        2512 => x"63662d15",
        2513 => x"8317c400",
        2514 => x"13f70748",
        2515 => x"63060708",
        2516 => x"83244401",
        2517 => x"83250401",
        2518 => x"832c0400",
        2519 => x"b3847403",
        2520 => x"b38cbc40",
        2521 => x"13871c00",
        2522 => x"3307a701",
        2523 => x"b3c48403",
        2524 => x"13860400",
        2525 => x"63f6e400",
        2526 => x"93040700",
        2527 => x"13060700",
        2528 => x"93f70740",
        2529 => x"6386070c",
        2530 => x"93050600",
        2531 => x"13050a00",
        2532 => x"eff0dfc0",
        2533 => x"13090500",
        2534 => x"630a050c",
        2535 => x"83250401",
        2536 => x"13860c00",
        2537 => x"efe09fc7",
        2538 => x"8357c400",
        2539 => x"93f7f7b7",
        2540 => x"93e70708",
        2541 => x"2316f400",
        2542 => x"23282401",
        2543 => x"232a9400",
        2544 => x"33099901",
        2545 => x"b3849441",
        2546 => x"23202401",
        2547 => x"23249400",
        2548 => x"13090d00",
        2549 => x"93040d00",
        2550 => x"03250400",
        2551 => x"13860400",
        2552 => x"93050b00",
        2553 => x"efe0dfc5",
        2554 => x"83278400",
        2555 => x"b3872741",
        2556 => x"2324f400",
        2557 => x"83270400",
        2558 => x"b3879700",
        2559 => x"2320f400",
        2560 => x"83a78900",
        2561 => x"b387a741",
        2562 => x"23a4f900",
        2563 => x"e39e07f0",
        2564 => x"13050000",
        2565 => x"8320c102",
        2566 => x"03248102",
        2567 => x"23a20900",
        2568 => x"83244102",
        2569 => x"03290102",
        2570 => x"8329c101",
        2571 => x"032a8101",
        2572 => x"832a4101",
        2573 => x"032b0101",
        2574 => x"832bc100",
        2575 => x"032c8100",
        2576 => x"832c4100",
        2577 => x"032d0100",
        2578 => x"13010103",
        2579 => x"67800000",
        2580 => x"13050a00",
        2581 => x"ef009041",
        2582 => x"13090500",
        2583 => x"e31e05f4",
        2584 => x"83250401",
        2585 => x"13050a00",
        2586 => x"eff09f9b",
        2587 => x"9307c000",
        2588 => x"2320fa00",
        2589 => x"8357c400",
        2590 => x"1305f0ff",
        2591 => x"93e70704",
        2592 => x"2316f400",
        2593 => x"23a40900",
        2594 => x"6ff0dff8",
        2595 => x"13090d00",
        2596 => x"6ff05ff4",
        2597 => x"83d7c500",
        2598 => x"130101f6",
        2599 => x"232c8108",
        2600 => x"232a9108",
        2601 => x"23282109",
        2602 => x"23244109",
        2603 => x"232e1108",
        2604 => x"23263109",
        2605 => x"23225109",
        2606 => x"23206109",
        2607 => x"232e7107",
        2608 => x"232c8107",
        2609 => x"232a9107",
        2610 => x"93f70708",
        2611 => x"130a0500",
        2612 => x"13890500",
        2613 => x"93040600",
        2614 => x"13840600",
        2615 => x"63840706",
        2616 => x"83a70501",
        2617 => x"63900706",
        2618 => x"93050004",
        2619 => x"eff01fab",
        2620 => x"2320a900",
        2621 => x"2328a900",
        2622 => x"63120504",
        2623 => x"9307c000",
        2624 => x"2320fa00",
        2625 => x"1305f0ff",
        2626 => x"8320c109",
        2627 => x"03248109",
        2628 => x"83244109",
        2629 => x"03290109",
        2630 => x"8329c108",
        2631 => x"032a8108",
        2632 => x"832a4108",
        2633 => x"032b0108",
        2634 => x"832bc107",
        2635 => x"032c8107",
        2636 => x"832c4107",
        2637 => x"1301010a",
        2638 => x"67800000",
        2639 => x"93070004",
        2640 => x"232af900",
        2641 => x"93070002",
        2642 => x"a304f102",
        2643 => x"93070003",
        2644 => x"23220102",
        2645 => x"2305f102",
        2646 => x"23268100",
        2647 => x"930b5002",
        2648 => x"930af0ff",
        2649 => x"130c1000",
        2650 => x"130ba000",
        2651 => x"13840400",
        2652 => x"83470400",
        2653 => x"63840700",
        2654 => x"6396770d",
        2655 => x"b30c9440",
        2656 => x"63049402",
        2657 => x"93860c00",
        2658 => x"13860400",
        2659 => x"93050900",
        2660 => x"13050a00",
        2661 => x"eff0dfbc",
        2662 => x"63045525",
        2663 => x"83274102",
        2664 => x"b3879701",
        2665 => x"2322f102",
        2666 => x"83470400",
        2667 => x"638a0722",
        2668 => x"93041400",
        2669 => x"23280100",
        2670 => x"232e0100",
        2671 => x"232a5101",
        2672 => x"232c0100",
        2673 => x"a3090104",
        2674 => x"23240106",
        2675 => x"b74c0000",
        2676 => x"83c50400",
        2677 => x"13065000",
        2678 => x"13858cbb",
        2679 => x"ef00901d",
        2680 => x"03270101",
        2681 => x"93070500",
        2682 => x"13841400",
        2683 => x"63100506",
        2684 => x"93770701",
        2685 => x"63860700",
        2686 => x"93070002",
        2687 => x"a309f104",
        2688 => x"93778700",
        2689 => x"63860700",
        2690 => x"9307b002",
        2691 => x"a309f104",
        2692 => x"83c60400",
        2693 => x"9307a002",
        2694 => x"6388f604",
        2695 => x"8327c101",
        2696 => x"13840400",
        2697 => x"93060000",
        2698 => x"13069000",
        2699 => x"03470400",
        2700 => x"93051400",
        2701 => x"130707fd",
        2702 => x"637ce608",
        2703 => x"63900604",
        2704 => x"6f004005",
        2705 => x"13041400",
        2706 => x"6ff09ff2",
        2707 => x"93868cbb",
        2708 => x"b387d740",
        2709 => x"b317fc00",
        2710 => x"b3e7e700",
        2711 => x"2328f100",
        2712 => x"93040400",
        2713 => x"6ff0dff6",
        2714 => x"8327c100",
        2715 => x"93864700",
        2716 => x"83a70700",
        2717 => x"2326d100",
        2718 => x"63c60700",
        2719 => x"232ef100",
        2720 => x"6f004001",
        2721 => x"b307f040",
        2722 => x"13672700",
        2723 => x"232ef100",
        2724 => x"2328e100",
        2725 => x"03470400",
        2726 => x"9307e002",
        2727 => x"6318f706",
        2728 => x"03471400",
        2729 => x"9307a002",
        2730 => x"631ef702",
        2731 => x"8327c100",
        2732 => x"13042400",
        2733 => x"13874700",
        2734 => x"83a70700",
        2735 => x"2326e100",
        2736 => x"63d40700",
        2737 => x"9307f0ff",
        2738 => x"232af100",
        2739 => x"6f000004",
        2740 => x"b3876703",
        2741 => x"13840500",
        2742 => x"93061000",
        2743 => x"b387e700",
        2744 => x"6ff0dff4",
        2745 => x"13041400",
        2746 => x"232a0100",
        2747 => x"93060000",
        2748 => x"93070000",
        2749 => x"13069000",
        2750 => x"03470400",
        2751 => x"93051400",
        2752 => x"130707fd",
        2753 => x"6378e608",
        2754 => x"e39006fc",
        2755 => x"83450400",
        2756 => x"b7440000",
        2757 => x"13063000",
        2758 => x"138504bc",
        2759 => x"ef009009",
        2760 => x"63020502",
        2761 => x"83270101",
        2762 => x"938404bc",
        2763 => x"33059540",
        2764 => x"13070004",
        2765 => x"3317a700",
        2766 => x"b3e7e700",
        2767 => x"13041400",
        2768 => x"2328f100",
        2769 => x"83450400",
        2770 => x"37450000",
        2771 => x"13066000",
        2772 => x"130545bc",
        2773 => x"93041400",
        2774 => x"2304b102",
        2775 => x"ef009005",
        2776 => x"630a0508",
        2777 => x"93070000",
        2778 => x"63980704",
        2779 => x"03270101",
        2780 => x"8327c100",
        2781 => x"13770710",
        2782 => x"63080702",
        2783 => x"93874700",
        2784 => x"2326f100",
        2785 => x"83274102",
        2786 => x"b3873701",
        2787 => x"2322f102",
        2788 => x"6ff0dfdd",
        2789 => x"b3876703",
        2790 => x"13840500",
        2791 => x"93061000",
        2792 => x"b387e700",
        2793 => x"6ff05ff5",
        2794 => x"93877700",
        2795 => x"93f787ff",
        2796 => x"93878700",
        2797 => x"6ff0dffc",
        2798 => x"b7260000",
        2799 => x"1307c100",
        2800 => x"93860656",
        2801 => x"13060900",
        2802 => x"93050101",
        2803 => x"13050a00",
        2804 => x"97000000",
        2805 => x"e7000000",
        2806 => x"93090500",
        2807 => x"e31455fb",
        2808 => x"8357c900",
        2809 => x"93f70704",
        2810 => x"e39e07d0",
        2811 => x"03254102",
        2812 => x"6ff09fd1",
        2813 => x"b7260000",
        2814 => x"1307c100",
        2815 => x"93860656",
        2816 => x"13060900",
        2817 => x"93050101",
        2818 => x"13050a00",
        2819 => x"ef00c01b",
        2820 => x"6ff09ffc",
        2821 => x"130101fd",
        2822 => x"232a5101",
        2823 => x"83a70501",
        2824 => x"930a0700",
        2825 => x"03a78500",
        2826 => x"23248102",
        2827 => x"23202103",
        2828 => x"232e3101",
        2829 => x"232c4101",
        2830 => x"23261102",
        2831 => x"23229102",
        2832 => x"23286101",
        2833 => x"23267101",
        2834 => x"93090500",
        2835 => x"13840500",
        2836 => x"13090600",
        2837 => x"138a0600",
        2838 => x"63d4e700",
        2839 => x"93070700",
        2840 => x"2320f900",
        2841 => x"03473404",
        2842 => x"63060700",
        2843 => x"93871700",
        2844 => x"2320f900",
        2845 => x"83270400",
        2846 => x"93f70702",
        2847 => x"63880700",
        2848 => x"83270900",
        2849 => x"93872700",
        2850 => x"2320f900",
        2851 => x"83240400",
        2852 => x"93f46400",
        2853 => x"639e0400",
        2854 => x"130b9401",
        2855 => x"930bf0ff",
        2856 => x"8327c400",
        2857 => x"03270900",
        2858 => x"b387e740",
        2859 => x"63c4f408",
        2860 => x"83473404",
        2861 => x"b336f000",
        2862 => x"83270400",
        2863 => x"93f70702",
        2864 => x"6392070c",
        2865 => x"13063404",
        2866 => x"93050a00",
        2867 => x"13850900",
        2868 => x"e7800a00",
        2869 => x"9307f0ff",
        2870 => x"630af506",
        2871 => x"83270400",
        2872 => x"13074000",
        2873 => x"93040000",
        2874 => x"93f76700",
        2875 => x"639ee700",
        2876 => x"83270900",
        2877 => x"8324c400",
        2878 => x"b384f440",
        2879 => x"93c7f4ff",
        2880 => x"93d7f741",
        2881 => x"b3f4f400",
        2882 => x"83278400",
        2883 => x"03270401",
        2884 => x"6356f700",
        2885 => x"b387e740",
        2886 => x"b384f400",
        2887 => x"13090000",
        2888 => x"1304a401",
        2889 => x"130bf0ff",
        2890 => x"63902409",
        2891 => x"13050000",
        2892 => x"6f000002",
        2893 => x"93061000",
        2894 => x"13060b00",
        2895 => x"93050a00",
        2896 => x"13850900",
        2897 => x"e7800a00",
        2898 => x"631a7503",
        2899 => x"1305f0ff",
        2900 => x"8320c102",
        2901 => x"03248102",
        2902 => x"83244102",
        2903 => x"03290102",
        2904 => x"8329c101",
        2905 => x"032a8101",
        2906 => x"832a4101",
        2907 => x"032b0101",
        2908 => x"832bc100",
        2909 => x"13010103",
        2910 => x"67800000",
        2911 => x"93841400",
        2912 => x"6ff01ff2",
        2913 => x"3307d400",
        2914 => x"13060003",
        2915 => x"a301c704",
        2916 => x"03475404",
        2917 => x"93871600",
        2918 => x"b307f400",
        2919 => x"93862600",
        2920 => x"a381e704",
        2921 => x"6ff01ff2",
        2922 => x"93061000",
        2923 => x"13060400",
        2924 => x"93050a00",
        2925 => x"13850900",
        2926 => x"e7800a00",
        2927 => x"e30865f9",
        2928 => x"13091900",
        2929 => x"6ff05ff6",
        2930 => x"130101fd",
        2931 => x"23248102",
        2932 => x"23229102",
        2933 => x"23202103",
        2934 => x"232e3101",
        2935 => x"23261102",
        2936 => x"232c4101",
        2937 => x"232a5101",
        2938 => x"23286101",
        2939 => x"83c88501",
        2940 => x"93078007",
        2941 => x"93040500",
        2942 => x"13840500",
        2943 => x"13090600",
        2944 => x"93890600",
        2945 => x"63ee1701",
        2946 => x"93072006",
        2947 => x"93863504",
        2948 => x"63ee1701",
        2949 => x"63840828",
        2950 => x"93078005",
        2951 => x"6380f822",
        2952 => x"930a2404",
        2953 => x"23011405",
        2954 => x"6f004004",
        2955 => x"9387d8f9",
        2956 => x"93f7f70f",
        2957 => x"13065001",
        2958 => x"e364f6fe",
        2959 => x"37460000",
        2960 => x"93972700",
        2961 => x"130646bf",
        2962 => x"b387c700",
        2963 => x"83a70700",
        2964 => x"67800700",
        2965 => x"83270700",
        2966 => x"938a2504",
        2967 => x"93864700",
        2968 => x"83a70700",
        2969 => x"2320d700",
        2970 => x"2381f504",
        2971 => x"93071000",
        2972 => x"6f008026",
        2973 => x"83a70500",
        2974 => x"03250700",
        2975 => x"13f60708",
        2976 => x"93054500",
        2977 => x"63060602",
        2978 => x"83270500",
        2979 => x"2320b700",
        2980 => x"37480000",
        2981 => x"63d80700",
        2982 => x"1307d002",
        2983 => x"b307f040",
        2984 => x"a301e404",
        2985 => x"1308c8bc",
        2986 => x"9308a000",
        2987 => x"6f004006",
        2988 => x"13f60704",
        2989 => x"83270500",
        2990 => x"2320b700",
        2991 => x"e30a06fc",
        2992 => x"93970701",
        2993 => x"93d70741",
        2994 => x"6ff09ffc",
        2995 => x"83a50500",
        2996 => x"03260700",
        2997 => x"13f50508",
        2998 => x"83270600",
        2999 => x"13064600",
        3000 => x"631a0500",
        3001 => x"93f50504",
        3002 => x"63860500",
        3003 => x"93970701",
        3004 => x"93d70701",
        3005 => x"2320c700",
        3006 => x"37480000",
        3007 => x"1307f006",
        3008 => x"1308c8bc",
        3009 => x"639ae814",
        3010 => x"93088000",
        3011 => x"a3010404",
        3012 => x"03274400",
        3013 => x"2324e400",
        3014 => x"634e0700",
        3015 => x"03260400",
        3016 => x"33e7e700",
        3017 => x"938a0600",
        3018 => x"1376b6ff",
        3019 => x"2320c400",
        3020 => x"63040702",
        3021 => x"938a0600",
        3022 => x"33f71703",
        3023 => x"938afaff",
        3024 => x"3307e800",
        3025 => x"03470700",
        3026 => x"2380ea00",
        3027 => x"13870700",
        3028 => x"b3d71703",
        3029 => x"e37217ff",
        3030 => x"93078000",
        3031 => x"6394f802",
        3032 => x"83270400",
        3033 => x"93f71700",
        3034 => x"638e0700",
        3035 => x"03274400",
        3036 => x"83270401",
        3037 => x"63c8e700",
        3038 => x"93070003",
        3039 => x"a38ffafe",
        3040 => x"938afaff",
        3041 => x"b3865641",
        3042 => x"2328d400",
        3043 => x"13870900",
        3044 => x"93060900",
        3045 => x"1306c100",
        3046 => x"93050400",
        3047 => x"13850400",
        3048 => x"eff05fc7",
        3049 => x"130af0ff",
        3050 => x"631e4513",
        3051 => x"1305f0ff",
        3052 => x"8320c102",
        3053 => x"03248102",
        3054 => x"83244102",
        3055 => x"03290102",
        3056 => x"8329c101",
        3057 => x"032a8101",
        3058 => x"832a4101",
        3059 => x"032b0101",
        3060 => x"13010103",
        3061 => x"67800000",
        3062 => x"83a70500",
        3063 => x"93e70702",
        3064 => x"23a0f500",
        3065 => x"37480000",
        3066 => x"93088007",
        3067 => x"130808be",
        3068 => x"a3021405",
        3069 => x"03260400",
        3070 => x"83250700",
        3071 => x"13750608",
        3072 => x"83a70500",
        3073 => x"93854500",
        3074 => x"631a0500",
        3075 => x"13750604",
        3076 => x"63060500",
        3077 => x"93970701",
        3078 => x"93d70701",
        3079 => x"2320b700",
        3080 => x"13771600",
        3081 => x"63060700",
        3082 => x"13660602",
        3083 => x"2320c400",
        3084 => x"638c0700",
        3085 => x"93080001",
        3086 => x"6ff05fed",
        3087 => x"37480000",
        3088 => x"1308c8bc",
        3089 => x"6ff0dffa",
        3090 => x"03270400",
        3091 => x"1377f7fd",
        3092 => x"2320e400",
        3093 => x"6ff01ffe",
        3094 => x"9308a000",
        3095 => x"6ff01feb",
        3096 => x"03a60500",
        3097 => x"83270700",
        3098 => x"83a54501",
        3099 => x"13780608",
        3100 => x"13854700",
        3101 => x"630a0800",
        3102 => x"2320a700",
        3103 => x"83a70700",
        3104 => x"23a0b700",
        3105 => x"6f008001",
        3106 => x"2320a700",
        3107 => x"13760604",
        3108 => x"83a70700",
        3109 => x"e30606fe",
        3110 => x"2390b700",
        3111 => x"23280400",
        3112 => x"938a0600",
        3113 => x"6ff09fee",
        3114 => x"83270700",
        3115 => x"03a64500",
        3116 => x"93050000",
        3117 => x"93864700",
        3118 => x"2320d700",
        3119 => x"83aa0700",
        3120 => x"13850a00",
        3121 => x"ef00002f",
        3122 => x"63060500",
        3123 => x"33055541",
        3124 => x"2322a400",
        3125 => x"83274400",
        3126 => x"2328f400",
        3127 => x"a3010404",
        3128 => x"6ff0dfea",
        3129 => x"83260401",
        3130 => x"13860a00",
        3131 => x"93050900",
        3132 => x"13850400",
        3133 => x"e7800900",
        3134 => x"e30a45eb",
        3135 => x"83270400",
        3136 => x"93f72700",
        3137 => x"63940704",
        3138 => x"8327c100",
        3139 => x"0325c400",
        3140 => x"e350f5ea",
        3141 => x"13850700",
        3142 => x"6ff09fe9",
        3143 => x"93061000",
        3144 => x"13060b00",
        3145 => x"93050900",
        3146 => x"13850400",
        3147 => x"e7800900",
        3148 => x"e30e45e7",
        3149 => x"938a1a00",
        3150 => x"8327c400",
        3151 => x"0327c100",
        3152 => x"b387e740",
        3153 => x"e3ccfafc",
        3154 => x"6ff01ffc",
        3155 => x"930a0000",
        3156 => x"130b9401",
        3157 => x"6ff05ffe",
        3158 => x"8397c500",
        3159 => x"130101fe",
        3160 => x"232c8100",
        3161 => x"232a9100",
        3162 => x"232e1100",
        3163 => x"23282101",
        3164 => x"23263101",
        3165 => x"13f78700",
        3166 => x"93040500",
        3167 => x"13840500",
        3168 => x"63120712",
        3169 => x"03a74500",
        3170 => x"6346e000",
        3171 => x"03a70504",
        3172 => x"6356e010",
        3173 => x"0327c402",
        3174 => x"63020710",
        3175 => x"03a90400",
        3176 => x"93963701",
        3177 => x"23a00400",
        3178 => x"63dc060a",
        3179 => x"03264405",
        3180 => x"8357c400",
        3181 => x"93f74700",
        3182 => x"638e0700",
        3183 => x"83274400",
        3184 => x"3306f640",
        3185 => x"83274403",
        3186 => x"63860700",
        3187 => x"83270404",
        3188 => x"3306f640",
        3189 => x"8327c402",
        3190 => x"83250402",
        3191 => x"93060000",
        3192 => x"13850400",
        3193 => x"e7800700",
        3194 => x"1307f0ff",
        3195 => x"8317c400",
        3196 => x"6312e502",
        3197 => x"83a60400",
        3198 => x"1307d001",
        3199 => x"636ad70e",
        3200 => x"37074020",
        3201 => x"13071700",
        3202 => x"3357d700",
        3203 => x"13771700",
        3204 => x"6300070e",
        3205 => x"03270401",
        3206 => x"23220400",
        3207 => x"2320e400",
        3208 => x"13973701",
        3209 => x"635c0700",
        3210 => x"9307f0ff",
        3211 => x"6316f500",
        3212 => x"83a70400",
        3213 => x"63940700",
        3214 => x"232aa404",
        3215 => x"83254403",
        3216 => x"23a02401",
        3217 => x"638c0504",
        3218 => x"93074404",
        3219 => x"6386f500",
        3220 => x"13850400",
        3221 => x"efe0dffc",
        3222 => x"232a0402",
        3223 => x"6f000004",
        3224 => x"83250402",
        3225 => x"13060000",
        3226 => x"93061000",
        3227 => x"13850400",
        3228 => x"e7000700",
        3229 => x"9307f0ff",
        3230 => x"13060500",
        3231 => x"e31af5f2",
        3232 => x"83a70400",
        3233 => x"e38607f2",
        3234 => x"1307d001",
        3235 => x"6386e700",
        3236 => x"13076001",
        3237 => x"639ce704",
        3238 => x"23a02401",
        3239 => x"13050000",
        3240 => x"6f00c005",
        3241 => x"83a90501",
        3242 => x"e38a09fe",
        3243 => x"03a90500",
        3244 => x"93f73700",
        3245 => x"23a03501",
        3246 => x"33093941",
        3247 => x"13070000",
        3248 => x"63940700",
        3249 => x"03a74501",
        3250 => x"2324e400",
        3251 => x"e35820fd",
        3252 => x"83278402",
        3253 => x"83250402",
        3254 => x"93060900",
        3255 => x"13860900",
        3256 => x"13850400",
        3257 => x"e7800700",
        3258 => x"6348a002",
        3259 => x"8317c400",
        3260 => x"93e70704",
        3261 => x"2316f400",
        3262 => x"1305f0ff",
        3263 => x"8320c101",
        3264 => x"03248101",
        3265 => x"83244101",
        3266 => x"03290101",
        3267 => x"8329c100",
        3268 => x"13010102",
        3269 => x"67800000",
        3270 => x"b389a900",
        3271 => x"3309a940",
        3272 => x"6ff0dffa",
        3273 => x"83a70501",
        3274 => x"638e0704",
        3275 => x"130101fe",
        3276 => x"232c8100",
        3277 => x"232e1100",
        3278 => x"13040500",
        3279 => x"630c0500",
        3280 => x"83270502",
        3281 => x"63980700",
        3282 => x"2326b100",
        3283 => x"efe05f85",
        3284 => x"8325c100",
        3285 => x"8397c500",
        3286 => x"638c0700",
        3287 => x"13050400",
        3288 => x"03248101",
        3289 => x"8320c101",
        3290 => x"13010102",
        3291 => x"6ff0dfde",
        3292 => x"8320c101",
        3293 => x"03248101",
        3294 => x"13050000",
        3295 => x"13010102",
        3296 => x"67800000",
        3297 => x"13050000",
        3298 => x"67800000",
        3299 => x"93050500",
        3300 => x"631e0500",
        3301 => x"b7350000",
        3302 => x"37050020",
        3303 => x"13868181",
        3304 => x"93854532",
        3305 => x"13054502",
        3306 => x"6fe0df84",
        3307 => x"03a50187",
        3308 => x"6ff05ff7",
        3309 => x"93f5f50f",
        3310 => x"3306c500",
        3311 => x"6316c500",
        3312 => x"13050000",
        3313 => x"67800000",
        3314 => x"83470500",
        3315 => x"e38cb7fe",
        3316 => x"13051500",
        3317 => x"6ff09ffe",
        3318 => x"130101ff",
        3319 => x"23248100",
        3320 => x"23229100",
        3321 => x"13040500",
        3322 => x"13850500",
        3323 => x"93050600",
        3324 => x"23261100",
        3325 => x"23ac0186",
        3326 => x"ef00801d",
        3327 => x"9307f0ff",
        3328 => x"6318f500",
        3329 => x"83a78187",
        3330 => x"63840700",
        3331 => x"2320f400",
        3332 => x"8320c100",
        3333 => x"03248100",
        3334 => x"83244100",
        3335 => x"13010101",
        3336 => x"67800000",
        3337 => x"130101ff",
        3338 => x"23248100",
        3339 => x"23229100",
        3340 => x"13040500",
        3341 => x"13850500",
        3342 => x"23261100",
        3343 => x"23ac0186",
        3344 => x"ef004028",
        3345 => x"9307f0ff",
        3346 => x"6318f500",
        3347 => x"83a78187",
        3348 => x"63840700",
        3349 => x"2320f400",
        3350 => x"8320c100",
        3351 => x"03248100",
        3352 => x"83244100",
        3353 => x"13010101",
        3354 => x"67800000",
        3355 => x"130101fe",
        3356 => x"232c8100",
        3357 => x"232e1100",
        3358 => x"232a9100",
        3359 => x"23282101",
        3360 => x"23263101",
        3361 => x"23244101",
        3362 => x"13040600",
        3363 => x"63940502",
        3364 => x"03248101",
        3365 => x"8320c101",
        3366 => x"83244101",
        3367 => x"03290101",
        3368 => x"8329c100",
        3369 => x"032a8100",
        3370 => x"93050600",
        3371 => x"13010102",
        3372 => x"6fe0dfee",
        3373 => x"63180602",
        3374 => x"efe09fd6",
        3375 => x"93040000",
        3376 => x"8320c101",
        3377 => x"03248101",
        3378 => x"03290101",
        3379 => x"8329c100",
        3380 => x"032a8100",
        3381 => x"13850400",
        3382 => x"83244101",
        3383 => x"13010102",
        3384 => x"67800000",
        3385 => x"130a0500",
        3386 => x"93840500",
        3387 => x"ef008005",
        3388 => x"13090500",
        3389 => x"63668500",
        3390 => x"93571500",
        3391 => x"e3e287fc",
        3392 => x"93050400",
        3393 => x"13050a00",
        3394 => x"efe05fe9",
        3395 => x"93090500",
        3396 => x"63160500",
        3397 => x"93840900",
        3398 => x"6ff09ffa",
        3399 => x"13060400",
        3400 => x"63748900",
        3401 => x"13060900",
        3402 => x"93850400",
        3403 => x"13850900",
        3404 => x"efd0dfee",
        3405 => x"93850400",
        3406 => x"13050a00",
        3407 => x"efe05fce",
        3408 => x"6ff05ffd",
        3409 => x"83a7c5ff",
        3410 => x"1385c7ff",
        3411 => x"63d80700",
        3412 => x"b385a500",
        3413 => x"83a70500",
        3414 => x"3305f500",
        3415 => x"67800000",
        3416 => x"130101ff",
        3417 => x"23261100",
        3418 => x"23248100",
        3419 => x"93089003",
        3420 => x"73000000",
        3421 => x"13040500",
        3422 => x"635a0500",
        3423 => x"33048040",
        3424 => x"efe0dfbe",
        3425 => x"23208500",
        3426 => x"1304f0ff",
        3427 => x"8320c100",
        3428 => x"13050400",
        3429 => x"03248100",
        3430 => x"13010101",
        3431 => x"67800000",
        3432 => x"9308d005",
        3433 => x"73000000",
        3434 => x"63520502",
        3435 => x"130101ff",
        3436 => x"23248100",
        3437 => x"13040500",
        3438 => x"23261100",
        3439 => x"33048040",
        3440 => x"efe0dfba",
        3441 => x"23208500",
        3442 => x"6f000000",
        3443 => x"6f000000",
        3444 => x"130101fe",
        3445 => x"232a9100",
        3446 => x"232e1100",
        3447 => x"93040500",
        3448 => x"232c8100",
        3449 => x"93083019",
        3450 => x"13050000",
        3451 => x"93050100",
        3452 => x"73000000",
        3453 => x"13040500",
        3454 => x"635a0500",
        3455 => x"33048040",
        3456 => x"efe0dfb6",
        3457 => x"23208500",
        3458 => x"1304f0ff",
        3459 => x"83274100",
        3460 => x"03270100",
        3461 => x"8320c101",
        3462 => x"23a2f400",
        3463 => x"83278100",
        3464 => x"23a0e400",
        3465 => x"1307803e",
        3466 => x"b3c7e702",
        3467 => x"13050400",
        3468 => x"03248101",
        3469 => x"23a4f400",
        3470 => x"83244101",
        3471 => x"13010102",
        3472 => x"67800000",
        3473 => x"130101ff",
        3474 => x"23261100",
        3475 => x"23248100",
        3476 => x"9308e003",
        3477 => x"73000000",
        3478 => x"13040500",
        3479 => x"635a0500",
        3480 => x"33048040",
        3481 => x"efe09fb0",
        3482 => x"23208500",
        3483 => x"1304f0ff",
        3484 => x"8320c100",
        3485 => x"13050400",
        3486 => x"03248100",
        3487 => x"13010101",
        3488 => x"67800000",
        3489 => x"130101ff",
        3490 => x"23261100",
        3491 => x"23248100",
        3492 => x"9308f003",
        3493 => x"73000000",
        3494 => x"13040500",
        3495 => x"635a0500",
        3496 => x"33048040",
        3497 => x"efe09fac",
        3498 => x"23208500",
        3499 => x"1304f0ff",
        3500 => x"8320c100",
        3501 => x"13050400",
        3502 => x"03248100",
        3503 => x"13010101",
        3504 => x"67800000",
        3505 => x"93070500",
        3506 => x"03a54188",
        3507 => x"130101ff",
        3508 => x"23261100",
        3509 => x"631a0502",
        3510 => x"9308600d",
        3511 => x"73000000",
        3512 => x"9306f0ff",
        3513 => x"6310d502",
        3514 => x"efe05fa8",
        3515 => x"9307c000",
        3516 => x"2320f500",
        3517 => x"1305f0ff",
        3518 => x"8320c100",
        3519 => x"13010101",
        3520 => x"67800000",
        3521 => x"23a2a188",
        3522 => x"9308600d",
        3523 => x"3385a700",
        3524 => x"73000000",
        3525 => x"93060500",
        3526 => x"03a54188",
        3527 => x"b387a700",
        3528 => x"e394f6fc",
        3529 => x"23a2d188",
        3530 => x"6ff01ffd",
        3531 => x"130101ff",
        3532 => x"23261100",
        3533 => x"23248100",
        3534 => x"93080004",
        3535 => x"73000000",
        3536 => x"13040500",
        3537 => x"635a0500",
        3538 => x"33048040",
        3539 => x"efe01fa2",
        3540 => x"23208500",
        3541 => x"1304f0ff",
        3542 => x"8320c100",
        3543 => x"13050400",
        3544 => x"03248100",
        3545 => x"13010101",
        3546 => x"67800000",
        3547 => x"10000000",
        3548 => x"00000000",
        3549 => x"037a5200",
        3550 => x"017c0101",
        3551 => x"1b0c0200",
        3552 => x"10000000",
        3553 => x"18000000",
        3554 => x"f8cfffff",
        3555 => x"74040000",
        3556 => x"00000000",
        3557 => x"10000000",
        3558 => x"00000000",
        3559 => x"037a5200",
        3560 => x"017c0101",
        3561 => x"1b0c0200",
        3562 => x"10000000",
        3563 => x"18000000",
        3564 => x"44d4ffff",
        3565 => x"2c040000",
        3566 => x"00000000",
        3567 => x"10000000",
        3568 => x"00000000",
        3569 => x"037a5200",
        3570 => x"017c0101",
        3571 => x"1b0c0200",
        3572 => x"10000000",
        3573 => x"18000000",
        3574 => x"48d8ffff",
        3575 => x"e0030000",
        3576 => x"00000000",
        3577 => x"30313233",
        3578 => x"34353637",
        3579 => x"38396162",
        3580 => x"63646566",
        3581 => x"00000000",
        3582 => x"a0040000",
        3583 => x"d8030000",
        3584 => x"d8030000",
        3585 => x"d8030000",
        3586 => x"ac040000",
        3587 => x"d8030000",
        3588 => x"d8030000",
        3589 => x"d8030000",
        3590 => x"d8030000",
        3591 => x"d8030000",
        3592 => x"d8030000",
        3593 => x"d8030000",
        3594 => x"d8030000",
        3595 => x"d8030000",
        3596 => x"d8030000",
        3597 => x"b8040000",
        3598 => x"d8030000",
        3599 => x"c4040000",
        3600 => x"d0040000",
        3601 => x"d8030000",
        3602 => x"dc040000",
        3603 => x"e8040000",
        3604 => x"d8030000",
        3605 => x"f4040000",
        3606 => x"94040000",
        3607 => x"d8030000",
        3608 => x"d8030000",
        3609 => x"d8030000",
        3610 => x"00050000",
        3611 => x"d8030000",
        3612 => x"d8030000",
        3613 => x"d8030000",
        3614 => x"d8030000",
        3615 => x"d8030000",
        3616 => x"d8030000",
        3617 => x"d8030000",
        3618 => x"10050000",
        3619 => x"a8050000",
        3620 => x"7c050000",
        3621 => x"7c050000",
        3622 => x"7c050000",
        3623 => x"7c050000",
        3624 => x"08060000",
        3625 => x"3c060000",
        3626 => x"14060000",
        3627 => x"7c050000",
        3628 => x"7c050000",
        3629 => x"7c050000",
        3630 => x"7c050000",
        3631 => x"7c050000",
        3632 => x"7c050000",
        3633 => x"7c050000",
        3634 => x"7c050000",
        3635 => x"7c050000",
        3636 => x"7c050000",
        3637 => x"7c050000",
        3638 => x"7c050000",
        3639 => x"7c050000",
        3640 => x"7c050000",
        3641 => x"94050000",
        3642 => x"94050000",
        3643 => x"7c050000",
        3644 => x"7c050000",
        3645 => x"7c050000",
        3646 => x"7c050000",
        3647 => x"7c050000",
        3648 => x"7c050000",
        3649 => x"7c050000",
        3650 => x"7c050000",
        3651 => x"7c050000",
        3652 => x"7c050000",
        3653 => x"7c050000",
        3654 => x"7c050000",
        3655 => x"08060000",
        3656 => x"a8050000",
        3657 => x"f0050000",
        3658 => x"d8050000",
        3659 => x"7c050000",
        3660 => x"7c050000",
        3661 => x"7c050000",
        3662 => x"7c050000",
        3663 => x"7c050000",
        3664 => x"7c050000",
        3665 => x"c0050000",
        3666 => x"7c050000",
        3667 => x"7c050000",
        3668 => x"7c050000",
        3669 => x"7c050000",
        3670 => x"94050000",
        3671 => x"94050000",
        3672 => x"00010202",
        3673 => x"03030303",
        3674 => x"04040404",
        3675 => x"04040404",
        3676 => x"05050505",
        3677 => x"05050505",
        3678 => x"05050505",
        3679 => x"05050505",
        3680 => x"06060606",
        3681 => x"06060606",
        3682 => x"06060606",
        3683 => x"06060606",
        3684 => x"06060606",
        3685 => x"06060606",
        3686 => x"06060606",
        3687 => x"06060606",
        3688 => x"07070707",
        3689 => x"07070707",
        3690 => x"07070707",
        3691 => x"07070707",
        3692 => x"07070707",
        3693 => x"07070707",
        3694 => x"07070707",
        3695 => x"07070707",
        3696 => x"07070707",
        3697 => x"07070707",
        3698 => x"07070707",
        3699 => x"07070707",
        3700 => x"07070707",
        3701 => x"07070707",
        3702 => x"07070707",
        3703 => x"07070707",
        3704 => x"08080808",
        3705 => x"08080808",
        3706 => x"08080808",
        3707 => x"08080808",
        3708 => x"08080808",
        3709 => x"08080808",
        3710 => x"08080808",
        3711 => x"08080808",
        3712 => x"08080808",
        3713 => x"08080808",
        3714 => x"08080808",
        3715 => x"08080808",
        3716 => x"08080808",
        3717 => x"08080808",
        3718 => x"08080808",
        3719 => x"08080808",
        3720 => x"08080808",
        3721 => x"08080808",
        3722 => x"08080808",
        3723 => x"08080808",
        3724 => x"08080808",
        3725 => x"08080808",
        3726 => x"08080808",
        3727 => x"08080808",
        3728 => x"08080808",
        3729 => x"08080808",
        3730 => x"08080808",
        3731 => x"08080808",
        3732 => x"08080808",
        3733 => x"08080808",
        3734 => x"08080808",
        3735 => x"08080808",
        3736 => x"0d0a4542",
        3737 => x"5245414b",
        3738 => x"21206d65",
        3739 => x"7063203d",
        3740 => x"20000000",
        3741 => x"20696e73",
        3742 => x"6e203d20",
        3743 => x"00000000",
        3744 => x"0d0a0000",
        3745 => x"0d0a0a44",
        3746 => x"6973706c",
        3747 => x"6179696e",
        3748 => x"67207468",
        3749 => x"65207469",
        3750 => x"6d652070",
        3751 => x"61737365",
        3752 => x"64207369",
        3753 => x"6e636520",
        3754 => x"72657365",
        3755 => x"740d0a0a",
        3756 => x"00000000",
        3757 => x"4f6e2d63",
        3758 => x"68697020",
        3759 => x"64656275",
        3760 => x"67676572",
        3761 => x"20666f75",
        3762 => x"6e642c20",
        3763 => x"736b6970",
        3764 => x"70696e67",
        3765 => x"20454252",
        3766 => x"45414b20",
        3767 => x"696e7374",
        3768 => x"72756374",
        3769 => x"696f6e0d",
        3770 => x"0a0d0a00",
        3771 => x"2530356c",
        3772 => x"643a2530",
        3773 => x"366c6420",
        3774 => x"20202530",
        3775 => x"326c643a",
        3776 => x"2530326c",
        3777 => x"643a2530",
        3778 => x"326c640d",
        3779 => x"00000000",
        3780 => x"696e7465",
        3781 => x"72727570",
        3782 => x"745f6469",
        3783 => x"72656374",
        3784 => x"00000000",
        3785 => x"54485541",
        3786 => x"53205249",
        3787 => x"53432d56",
        3788 => x"20525633",
        3789 => x"32494d20",
        3790 => x"62617265",
        3791 => x"206d6574",
        3792 => x"616c2070",
        3793 => x"726f6365",
        3794 => x"73736f72",
        3795 => x"00000000",
        3796 => x"54686520",
        3797 => x"48616775",
        3798 => x"6520556e",
        3799 => x"69766572",
        3800 => x"73697479",
        3801 => x"206f6620",
        3802 => x"4170706c",
        3803 => x"69656420",
        3804 => x"53636965",
        3805 => x"6e636573",
        3806 => x"00000000",
        3807 => x"44657061",
        3808 => x"72746d65",
        3809 => x"6e74206f",
        3810 => x"6620456c",
        3811 => x"65637472",
        3812 => x"6963616c",
        3813 => x"20456e67",
        3814 => x"696e6565",
        3815 => x"72696e67",
        3816 => x"00000000",
        3817 => x"4a2e452e",
        3818 => x"4a2e206f",
        3819 => x"70206465",
        3820 => x"6e204272",
        3821 => x"6f757700",
        3822 => x"232d302b",
        3823 => x"20000000",
        3824 => x"686c4c00",
        3825 => x"65666745",
        3826 => x"46470000",
        3827 => x"30313233",
        3828 => x"34353637",
        3829 => x"38394142",
        3830 => x"43444546",
        3831 => x"00000000",
        3832 => x"30313233",
        3833 => x"34353637",
        3834 => x"38396162",
        3835 => x"63646566",
        3836 => x"00000000",
        3837 => x"542e0000",
        3838 => x"742e0000",
        3839 => x"202e0000",
        3840 => x"202e0000",
        3841 => x"202e0000",
        3842 => x"202e0000",
        3843 => x"742e0000",
        3844 => x"202e0000",
        3845 => x"202e0000",
        3846 => x"202e0000",
        3847 => x"202e0000",
        3848 => x"60300000",
        3849 => x"cc2e0000",
        3850 => x"d82f0000",
        3851 => x"202e0000",
        3852 => x"202e0000",
        3853 => x"a8300000",
        3854 => x"202e0000",
        3855 => x"cc2e0000",
        3856 => x"202e0000",
        3857 => x"202e0000",
        3858 => x"e42f0000",
        3859 => x"103b0000",
        3860 => x"243b0000",
        3861 => x"503b0000",
        3862 => x"7c3b0000",
        3863 => x"a43b0000",
        3864 => x"00000000",
        3865 => x"00000000",
        3866 => x"03000000",
        3867 => x"88000020",
        3868 => x"00000000",
        3869 => x"88000020",
        3870 => x"f0000020",
        3871 => x"58010020",
        3872 => x"00000000",
        3873 => x"00000000",
        3874 => x"00000000",
        3875 => x"00000000",
        3876 => x"00000000",
        3877 => x"00000000",
        3878 => x"00000000",
        3879 => x"00000000",
        3880 => x"00000000",
        3881 => x"00000000",
        3882 => x"00000000",
        3883 => x"00000000",
        3884 => x"00000000",
        3885 => x"00000000",
        3886 => x"00000000",
        3887 => x"24000020",
        3888 => x"00000000"
            );
end package rom_image;
