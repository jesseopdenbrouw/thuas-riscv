-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Sat Nov 23 16:00:52 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382c22e",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"13060500",
           9 => x"93878186",
          10 => x"637cf600",
          11 => x"b7350000",
          12 => x"3386c740",
          13 => x"13050500",
          14 => x"938585e5",
          15 => x"ef108035",
          16 => x"13868186",
          17 => x"9387419b",
          18 => x"637af600",
          19 => x"3386c740",
          20 => x"13858186",
          21 => x"93050000",
          22 => x"ef100032",
          23 => x"ef10501c",
          24 => x"b7050020",
          25 => x"93850500",
          26 => x"13060000",
          27 => x"13055000",
          28 => x"ef10c052",
          29 => x"ef10900f",
          30 => x"6f104047",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef10804b",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"b7370000",
          40 => x"232c4101",
          41 => x"130a0500",
          42 => x"1385c7c6",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"37390000",
          50 => x"ef104049",
          51 => x"13044100",
          52 => x"93070400",
          53 => x"9309c1ff",
          54 => x"1309099f",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef10c045",
          65 => x"37350000",
          66 => x"130505c8",
          67 => x"ef100045",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef108042",
          78 => x"37350000",
          79 => x"1305c5c8",
          80 => x"ef10c041",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74760",
          91 => x"93860700",
          92 => x"1377f7fe",
          93 => x"23a2e760",
          94 => x"83a74700",
          95 => x"93c71700",
          96 => x"23a2f600",
          97 => x"67800000",
          98 => x"370700f0",
          99 => x"83274700",
         100 => x"93e70720",
         101 => x"2322f700",
         102 => x"6f000000",
         103 => x"b71700f0",
         104 => x"93850700",
         105 => x"938505a0",
         106 => x"938747a0",
         107 => x"83a60700",
         108 => x"03a60500",
         109 => x"03a70700",
         110 => x"e31ad7fe",
         111 => x"b7870100",
         112 => x"b71600f0",
         113 => x"1305f0ff",
         114 => x"9387076a",
         115 => x"23a6a6a0",
         116 => x"b307f600",
         117 => x"23a4a6a0",
         118 => x"33b6c700",
         119 => x"23a4f6a0",
         120 => x"3306e600",
         121 => x"23a6c6a0",
         122 => x"370700f0",
         123 => x"83274700",
         124 => x"93c72700",
         125 => x"2322f700",
         126 => x"67800000",
         127 => x"b70700f0",
         128 => x"03a74710",
         129 => x"b70600f0",
         130 => x"93870710",
         131 => x"13778700",
         132 => x"630a0700",
         133 => x"03a74600",
         134 => x"13478700",
         135 => x"23a2e600",
         136 => x"83a78700",
         137 => x"67800000",
         138 => x"b70700f0",
         139 => x"03a74770",
         140 => x"93860700",
         141 => x"1377f7f0",
         142 => x"23a2e770",
         143 => x"83a74700",
         144 => x"93c74700",
         145 => x"23a2f600",
         146 => x"67800000",
         147 => x"b70700f0",
         148 => x"03a74740",
         149 => x"93860700",
         150 => x"137777ff",
         151 => x"23a2e740",
         152 => x"83a74700",
         153 => x"93c70701",
         154 => x"23a2f600",
         155 => x"67800000",
         156 => x"b70700f0",
         157 => x"03a74720",
         158 => x"93860700",
         159 => x"137777ff",
         160 => x"23a2e720",
         161 => x"83a74700",
         162 => x"93c70702",
         163 => x"23a2f600",
         164 => x"67800000",
         165 => x"b70700f0",
         166 => x"03a74730",
         167 => x"93860700",
         168 => x"137777ff",
         169 => x"23a2e730",
         170 => x"83a74700",
         171 => x"93c70708",
         172 => x"23a2f600",
         173 => x"67800000",
         174 => x"b70700f0",
         175 => x"23ae0700",
         176 => x"03a74700",
         177 => x"13470704",
         178 => x"23a2e700",
         179 => x"67800000",
         180 => x"b71700f0",
         181 => x"23a00790",
         182 => x"370700f0",
         183 => x"83274700",
         184 => x"93c70710",
         185 => x"2322f700",
         186 => x"67800000",
         187 => x"6f000000",
         188 => x"13050000",
         189 => x"67800000",
         190 => x"13050000",
         191 => x"67800000",
         192 => x"130101f7",
         193 => x"23221100",
         194 => x"23242100",
         195 => x"23263100",
         196 => x"23284100",
         197 => x"232a5100",
         198 => x"232c6100",
         199 => x"232e7100",
         200 => x"23208102",
         201 => x"23229102",
         202 => x"2324a102",
         203 => x"2326b102",
         204 => x"2328c102",
         205 => x"232ad102",
         206 => x"232ce102",
         207 => x"232ef102",
         208 => x"23200105",
         209 => x"23221105",
         210 => x"23242105",
         211 => x"23263105",
         212 => x"23284105",
         213 => x"232a5105",
         214 => x"232c6105",
         215 => x"232e7105",
         216 => x"23208107",
         217 => x"23229107",
         218 => x"2324a107",
         219 => x"2326b107",
         220 => x"2328c107",
         221 => x"232ad107",
         222 => x"232ce107",
         223 => x"232ef107",
         224 => x"f3222034",
         225 => x"23205108",
         226 => x"f3221034",
         227 => x"23225108",
         228 => x"83a20200",
         229 => x"23245108",
         230 => x"f3223034",
         231 => x"23265108",
         232 => x"f3272034",
         233 => x"1307b000",
         234 => x"6374f70c",
         235 => x"37070080",
         236 => x"1307d7ff",
         237 => x"b387e700",
         238 => x"13078001",
         239 => x"636ef700",
         240 => x"37370000",
         241 => x"93972700",
         242 => x"130747a0",
         243 => x"b387e700",
         244 => x"83a70700",
         245 => x"67800700",
         246 => x"03258102",
         247 => x"83220108",
         248 => x"63c80200",
         249 => x"f3221034",
         250 => x"93824200",
         251 => x"73901234",
         252 => x"832fc107",
         253 => x"032f8107",
         254 => x"832e4107",
         255 => x"032e0107",
         256 => x"832dc106",
         257 => x"032d8106",
         258 => x"832c4106",
         259 => x"032c0106",
         260 => x"832bc105",
         261 => x"032b8105",
         262 => x"832a4105",
         263 => x"032a0105",
         264 => x"8329c104",
         265 => x"03298104",
         266 => x"83284104",
         267 => x"03280104",
         268 => x"8327c103",
         269 => x"03278103",
         270 => x"83264103",
         271 => x"03260103",
         272 => x"8325c102",
         273 => x"83244102",
         274 => x"03240102",
         275 => x"8323c101",
         276 => x"03238101",
         277 => x"83224101",
         278 => x"03220101",
         279 => x"8321c100",
         280 => x"03218100",
         281 => x"83204100",
         282 => x"13010109",
         283 => x"73002030",
         284 => x"93061000",
         285 => x"e3f2f6f6",
         286 => x"e360f7f6",
         287 => x"37370000",
         288 => x"93972700",
         289 => x"130787a6",
         290 => x"b387e700",
         291 => x"83a70700",
         292 => x"67800700",
         293 => x"eff09fdb",
         294 => x"03258102",
         295 => x"6ff01ff4",
         296 => x"eff01fe3",
         297 => x"03258102",
         298 => x"6ff05ff3",
         299 => x"eff01fcf",
         300 => x"03258102",
         301 => x"6ff09ff2",
         302 => x"eff01fe0",
         303 => x"03258102",
         304 => x"6ff0dff1",
         305 => x"eff01fca",
         306 => x"03258102",
         307 => x"6ff01ff1",
         308 => x"eff09fd5",
         309 => x"03258102",
         310 => x"6ff05ff0",
         311 => x"eff01fd2",
         312 => x"03258102",
         313 => x"6ff09fef",
         314 => x"eff0dfda",
         315 => x"03258102",
         316 => x"6ff0dfee",
         317 => x"eff0dfd7",
         318 => x"03258102",
         319 => x"6ff01fee",
         320 => x"13050100",
         321 => x"eff05fb9",
         322 => x"03258102",
         323 => x"6ff01fed",
         324 => x"9307900a",
         325 => x"6380f814",
         326 => x"63d81703",
         327 => x"9307600d",
         328 => x"638ef818",
         329 => x"938808c0",
         330 => x"9307f000",
         331 => x"63e01705",
         332 => x"b7370000",
         333 => x"938787a9",
         334 => x"93982800",
         335 => x"b388f800",
         336 => x"83a70800",
         337 => x"67800700",
         338 => x"938878fc",
         339 => x"93074002",
         340 => x"63ee1701",
         341 => x"b7370000",
         342 => x"938787ad",
         343 => x"93982800",
         344 => x"b388f800",
         345 => x"83a70800",
         346 => x"67800700",
         347 => x"ef10c04a",
         348 => x"93078005",
         349 => x"2320f500",
         350 => x"9307f0ff",
         351 => x"13850700",
         352 => x"6ff0dfe5",
         353 => x"b7270000",
         354 => x"23a2f500",
         355 => x"93070000",
         356 => x"13850700",
         357 => x"6ff09fe4",
         358 => x"93070000",
         359 => x"13850700",
         360 => x"6ff0dfe3",
         361 => x"ef104047",
         362 => x"93079000",
         363 => x"2320f500",
         364 => x"9307f0ff",
         365 => x"13850700",
         366 => x"6ff05fe2",
         367 => x"ef10c045",
         368 => x"9307f001",
         369 => x"2320f500",
         370 => x"9307f0ff",
         371 => x"13850700",
         372 => x"6ff0dfe0",
         373 => x"ef104044",
         374 => x"9307d000",
         375 => x"2320f500",
         376 => x"9307f0ff",
         377 => x"13850700",
         378 => x"6ff05fdf",
         379 => x"ef10c042",
         380 => x"93072000",
         381 => x"2320f500",
         382 => x"9307f0ff",
         383 => x"13850700",
         384 => x"6ff0dfdd",
         385 => x"13090600",
         386 => x"13840500",
         387 => x"635cc000",
         388 => x"b384c500",
         389 => x"eff05fa6",
         390 => x"2300a400",
         391 => x"13041400",
         392 => x"e39a84fe",
         393 => x"13050900",
         394 => x"6ff05fdb",
         395 => x"13090600",
         396 => x"13840500",
         397 => x"e358c0fe",
         398 => x"b384c500",
         399 => x"03450400",
         400 => x"13041400",
         401 => x"eff09fa3",
         402 => x"e39a84fe",
         403 => x"13050900",
         404 => x"6ff0dfd8",
         405 => x"13090000",
         406 => x"93040500",
         407 => x"13040900",
         408 => x"93090900",
         409 => x"93070900",
         410 => x"732410c8",
         411 => x"f32910c0",
         412 => x"f32710c8",
         413 => x"e31af4fe",
         414 => x"37460f00",
         415 => x"13060624",
         416 => x"93060000",
         417 => x"13850900",
         418 => x"93050400",
         419 => x"ef00d010",
         420 => x"37460f00",
         421 => x"23a4a400",
         422 => x"93050400",
         423 => x"13850900",
         424 => x"13060624",
         425 => x"93060000",
         426 => x"ef00404c",
         427 => x"23a0a400",
         428 => x"23a2b400",
         429 => x"13050900",
         430 => x"6ff05fd2",
         431 => x"63180500",
         432 => x"1385819b",
         433 => x"13050500",
         434 => x"6ff05fd1",
         435 => x"b7870020",
         436 => x"93870700",
         437 => x"13070040",
         438 => x"b387e740",
         439 => x"e364f5fe",
         440 => x"ef108033",
         441 => x"9307c000",
         442 => x"2320f500",
         443 => x"1305f0ff",
         444 => x"13050500",
         445 => x"6ff09fce",
         446 => x"13030500",
         447 => x"138e0500",
         448 => x"93080000",
         449 => x"63dc0500",
         450 => x"b337a000",
         451 => x"3307b040",
         452 => x"330ef740",
         453 => x"3303a040",
         454 => x"9308f0ff",
         455 => x"63dc0600",
         456 => x"b337c000",
         457 => x"b306d040",
         458 => x"93c8f8ff",
         459 => x"b386f640",
         460 => x"3306c040",
         461 => x"13070600",
         462 => x"13080300",
         463 => x"93070e00",
         464 => x"639c0628",
         465 => x"b7350000",
         466 => x"9385c5b6",
         467 => x"6376ce0e",
         468 => x"b7060100",
         469 => x"6378d60c",
         470 => x"93360610",
         471 => x"93b61600",
         472 => x"93963600",
         473 => x"3355d600",
         474 => x"b385a500",
         475 => x"83c50500",
         476 => x"13050002",
         477 => x"b386d500",
         478 => x"b305d540",
         479 => x"630cd500",
         480 => x"b317be00",
         481 => x"b356d300",
         482 => x"3317b600",
         483 => x"b3e7f600",
         484 => x"3318b300",
         485 => x"93550701",
         486 => x"33deb702",
         487 => x"13160701",
         488 => x"13560601",
         489 => x"b3f7b702",
         490 => x"13050e00",
         491 => x"3303c603",
         492 => x"93960701",
         493 => x"93570801",
         494 => x"b3e7d700",
         495 => x"63fe6700",
         496 => x"b307f700",
         497 => x"1305feff",
         498 => x"63e8e700",
         499 => x"63f66700",
         500 => x"1305eeff",
         501 => x"b387e700",
         502 => x"b3876740",
         503 => x"33d3b702",
         504 => x"13180801",
         505 => x"13580801",
         506 => x"b3f7b702",
         507 => x"b3066602",
         508 => x"93970701",
         509 => x"3368f800",
         510 => x"93070300",
         511 => x"637cd800",
         512 => x"33080701",
         513 => x"9307f3ff",
         514 => x"6366e800",
         515 => x"6374d800",
         516 => x"9307e3ff",
         517 => x"13150501",
         518 => x"3365f500",
         519 => x"93050000",
         520 => x"6f00000e",
         521 => x"37050001",
         522 => x"93068001",
         523 => x"e37ca6f2",
         524 => x"93060001",
         525 => x"6ff01ff3",
         526 => x"93060000",
         527 => x"630c0600",
         528 => x"b7070100",
         529 => x"637af60c",
         530 => x"93360610",
         531 => x"93b61600",
         532 => x"93963600",
         533 => x"b357d600",
         534 => x"b385f500",
         535 => x"83c70500",
         536 => x"b387d700",
         537 => x"93060002",
         538 => x"b385f640",
         539 => x"6390f60c",
         540 => x"b307ce40",
         541 => x"93051000",
         542 => x"13530701",
         543 => x"b3de6702",
         544 => x"13160701",
         545 => x"13560601",
         546 => x"93560801",
         547 => x"b3f76702",
         548 => x"13850e00",
         549 => x"330ed603",
         550 => x"93970701",
         551 => x"b3e7f600",
         552 => x"63fec701",
         553 => x"b307f700",
         554 => x"1385feff",
         555 => x"63e8e700",
         556 => x"63f6c701",
         557 => x"1385eeff",
         558 => x"b387e700",
         559 => x"b387c741",
         560 => x"33de6702",
         561 => x"13180801",
         562 => x"13580801",
         563 => x"b3f76702",
         564 => x"b306c603",
         565 => x"93970701",
         566 => x"3368f800",
         567 => x"93070e00",
         568 => x"637cd800",
         569 => x"33080701",
         570 => x"9307feff",
         571 => x"6366e800",
         572 => x"6374d800",
         573 => x"9307eeff",
         574 => x"13150501",
         575 => x"3365f500",
         576 => x"638a0800",
         577 => x"b337a000",
         578 => x"b305b040",
         579 => x"b385f540",
         580 => x"3305a040",
         581 => x"67800000",
         582 => x"b7070001",
         583 => x"93068001",
         584 => x"e37af6f2",
         585 => x"93060001",
         586 => x"6ff0dff2",
         587 => x"3317b600",
         588 => x"b356fe00",
         589 => x"13550701",
         590 => x"331ebe00",
         591 => x"b357f300",
         592 => x"b3e7c701",
         593 => x"33dea602",
         594 => x"13160701",
         595 => x"13560601",
         596 => x"3318b300",
         597 => x"b3f6a602",
         598 => x"3303c603",
         599 => x"93950601",
         600 => x"93d60701",
         601 => x"b3e6b600",
         602 => x"93050e00",
         603 => x"63fe6600",
         604 => x"b306d700",
         605 => x"9305feff",
         606 => x"63e8e600",
         607 => x"63f66600",
         608 => x"9305eeff",
         609 => x"b386e600",
         610 => x"b3866640",
         611 => x"33d3a602",
         612 => x"93970701",
         613 => x"93d70701",
         614 => x"b3f6a602",
         615 => x"33066602",
         616 => x"93960601",
         617 => x"b3e7d700",
         618 => x"93060300",
         619 => x"63fec700",
         620 => x"b307f700",
         621 => x"9306f3ff",
         622 => x"63e8e700",
         623 => x"63f6c700",
         624 => x"9306e3ff",
         625 => x"b387e700",
         626 => x"93950501",
         627 => x"b387c740",
         628 => x"b3e5d500",
         629 => x"6ff05fea",
         630 => x"6364de18",
         631 => x"b7070100",
         632 => x"63f4f604",
         633 => x"13b70610",
         634 => x"13371700",
         635 => x"13173700",
         636 => x"b7370000",
         637 => x"b3d5e600",
         638 => x"9387c7b6",
         639 => x"b387b700",
         640 => x"83c70700",
         641 => x"b387e700",
         642 => x"13070002",
         643 => x"b305f740",
         644 => x"6316f702",
         645 => x"13051000",
         646 => x"e3e4c6ef",
         647 => x"3335c300",
         648 => x"13351500",
         649 => x"6ff0dfed",
         650 => x"b7070001",
         651 => x"13078001",
         652 => x"e3f0f6fc",
         653 => x"13070001",
         654 => x"6ff09ffb",
         655 => x"3358f600",
         656 => x"b396b600",
         657 => x"3368d800",
         658 => x"3355fe00",
         659 => x"3317be00",
         660 => x"135e0801",
         661 => x"335fc503",
         662 => x"93160801",
         663 => x"93d60601",
         664 => x"b357f300",
         665 => x"b3e7e700",
         666 => x"13d70701",
         667 => x"3316b600",
         668 => x"3375c503",
         669 => x"b38ee603",
         670 => x"13150501",
         671 => x"3367a700",
         672 => x"13050f00",
         673 => x"637ed701",
         674 => x"3307e800",
         675 => x"1305ffff",
         676 => x"63680701",
         677 => x"6376d701",
         678 => x"1305efff",
         679 => x"33070701",
         680 => x"3307d741",
         681 => x"b35ec703",
         682 => x"93970701",
         683 => x"93d70701",
         684 => x"3377c703",
         685 => x"b386d603",
         686 => x"13170701",
         687 => x"b3e7e700",
         688 => x"13870e00",
         689 => x"63fed700",
         690 => x"b307f800",
         691 => x"1387feff",
         692 => x"63e80701",
         693 => x"63f6d700",
         694 => x"1387eeff",
         695 => x"b3870701",
         696 => x"13150501",
         697 => x"3365e500",
         698 => x"131e0601",
         699 => x"13170701",
         700 => x"13570701",
         701 => x"13580501",
         702 => x"135e0e01",
         703 => x"13560601",
         704 => x"b30ec703",
         705 => x"b387d740",
         706 => x"330ec803",
         707 => x"93d60e01",
         708 => x"3307c702",
         709 => x"3307c701",
         710 => x"3387e600",
         711 => x"3308c802",
         712 => x"6376c701",
         713 => x"b7060100",
         714 => x"3308d800",
         715 => x"93560701",
         716 => x"b3860601",
         717 => x"63e2d702",
         718 => x"e392d7ce",
         719 => x"939e0e01",
         720 => x"13170701",
         721 => x"93de0e01",
         722 => x"3313b300",
         723 => x"3307d701",
         724 => x"93050000",
         725 => x"e376e3da",
         726 => x"1305f5ff",
         727 => x"6ff01fcc",
         728 => x"93050000",
         729 => x"13050000",
         730 => x"6ff09fd9",
         731 => x"93080500",
         732 => x"13830500",
         733 => x"13070600",
         734 => x"13080500",
         735 => x"93870500",
         736 => x"63920628",
         737 => x"b7350000",
         738 => x"9385c5b6",
         739 => x"6376c30e",
         740 => x"b7060100",
         741 => x"6378d60c",
         742 => x"93360610",
         743 => x"93b61600",
         744 => x"93963600",
         745 => x"3355d600",
         746 => x"b385a500",
         747 => x"83c50500",
         748 => x"13050002",
         749 => x"b386d500",
         750 => x"b305d540",
         751 => x"630cd500",
         752 => x"b317b300",
         753 => x"b3d6d800",
         754 => x"3317b600",
         755 => x"b3e7f600",
         756 => x"3398b800",
         757 => x"93550701",
         758 => x"33d3b702",
         759 => x"13160701",
         760 => x"13560601",
         761 => x"b3f7b702",
         762 => x"13050300",
         763 => x"b3086602",
         764 => x"93960701",
         765 => x"93570801",
         766 => x"b3e7d700",
         767 => x"63fe1701",
         768 => x"b307f700",
         769 => x"1305f3ff",
         770 => x"63e8e700",
         771 => x"63f61701",
         772 => x"1305e3ff",
         773 => x"b387e700",
         774 => x"b3871741",
         775 => x"b3d8b702",
         776 => x"13180801",
         777 => x"13580801",
         778 => x"b3f7b702",
         779 => x"b3061603",
         780 => x"93970701",
         781 => x"3368f800",
         782 => x"93870800",
         783 => x"637cd800",
         784 => x"33080701",
         785 => x"9387f8ff",
         786 => x"6366e800",
         787 => x"6374d800",
         788 => x"9387e8ff",
         789 => x"13150501",
         790 => x"3365f500",
         791 => x"93050000",
         792 => x"67800000",
         793 => x"37050001",
         794 => x"93068001",
         795 => x"e37ca6f2",
         796 => x"93060001",
         797 => x"6ff01ff3",
         798 => x"93060000",
         799 => x"630c0600",
         800 => x"b7070100",
         801 => x"6370f60c",
         802 => x"93360610",
         803 => x"93b61600",
         804 => x"93963600",
         805 => x"b357d600",
         806 => x"b385f500",
         807 => x"83c70500",
         808 => x"b387d700",
         809 => x"93060002",
         810 => x"b385f640",
         811 => x"6396f60a",
         812 => x"b307c340",
         813 => x"93051000",
         814 => x"93580701",
         815 => x"33de1703",
         816 => x"13160701",
         817 => x"13560601",
         818 => x"93560801",
         819 => x"b3f71703",
         820 => x"13050e00",
         821 => x"3303c603",
         822 => x"93970701",
         823 => x"b3e7f600",
         824 => x"63fe6700",
         825 => x"b307f700",
         826 => x"1305feff",
         827 => x"63e8e700",
         828 => x"63f66700",
         829 => x"1305eeff",
         830 => x"b387e700",
         831 => x"b3876740",
         832 => x"33d31703",
         833 => x"13180801",
         834 => x"13580801",
         835 => x"b3f71703",
         836 => x"b3066602",
         837 => x"93970701",
         838 => x"3368f800",
         839 => x"93070300",
         840 => x"637cd800",
         841 => x"33080701",
         842 => x"9307f3ff",
         843 => x"6366e800",
         844 => x"6374d800",
         845 => x"9307e3ff",
         846 => x"13150501",
         847 => x"3365f500",
         848 => x"67800000",
         849 => x"b7070001",
         850 => x"93068001",
         851 => x"e374f6f4",
         852 => x"93060001",
         853 => x"6ff01ff4",
         854 => x"3317b600",
         855 => x"b356f300",
         856 => x"13550701",
         857 => x"3313b300",
         858 => x"b3d7f800",
         859 => x"b3e76700",
         860 => x"33d3a602",
         861 => x"13160701",
         862 => x"13560601",
         863 => x"3398b800",
         864 => x"b3f6a602",
         865 => x"b3086602",
         866 => x"93950601",
         867 => x"93d60701",
         868 => x"b3e6b600",
         869 => x"93050300",
         870 => x"63fe1601",
         871 => x"b306d700",
         872 => x"9305f3ff",
         873 => x"63e8e600",
         874 => x"63f61601",
         875 => x"9305e3ff",
         876 => x"b386e600",
         877 => x"b3861641",
         878 => x"b3d8a602",
         879 => x"93970701",
         880 => x"93d70701",
         881 => x"b3f6a602",
         882 => x"33061603",
         883 => x"93960601",
         884 => x"b3e7d700",
         885 => x"93860800",
         886 => x"63fec700",
         887 => x"b307f700",
         888 => x"9386f8ff",
         889 => x"63e8e700",
         890 => x"63f6c700",
         891 => x"9386e8ff",
         892 => x"b387e700",
         893 => x"93950501",
         894 => x"b387c740",
         895 => x"b3e5d500",
         896 => x"6ff09feb",
         897 => x"63e4d518",
         898 => x"b7070100",
         899 => x"63f4f604",
         900 => x"93b70610",
         901 => x"93b71700",
         902 => x"93973700",
         903 => x"37370000",
         904 => x"b3d5f600",
         905 => x"1307c7b6",
         906 => x"3307b700",
         907 => x"03470700",
         908 => x"3307f700",
         909 => x"93070002",
         910 => x"b385e740",
         911 => x"6396e702",
         912 => x"13051000",
         913 => x"e3ee66e0",
         914 => x"33b5c800",
         915 => x"13351500",
         916 => x"67800000",
         917 => x"37070001",
         918 => x"93078001",
         919 => x"e3f0e6fc",
         920 => x"93070001",
         921 => x"6ff09ffb",
         922 => x"3355e600",
         923 => x"b396b600",
         924 => x"b357e300",
         925 => x"3365d500",
         926 => x"3313b300",
         927 => x"33d7e800",
         928 => x"33676700",
         929 => x"13530501",
         930 => x"b3de6702",
         931 => x"13180501",
         932 => x"13580801",
         933 => x"93560701",
         934 => x"3316b600",
         935 => x"b3f76702",
         936 => x"330ed803",
         937 => x"93970701",
         938 => x"b3e6f600",
         939 => x"93870e00",
         940 => x"63fec601",
         941 => x"b306d500",
         942 => x"9387feff",
         943 => x"63e8a600",
         944 => x"63f6c601",
         945 => x"9387eeff",
         946 => x"b386a600",
         947 => x"b386c641",
         948 => x"33de6602",
         949 => x"13170701",
         950 => x"13570701",
         951 => x"b3f66602",
         952 => x"3308c803",
         953 => x"93960601",
         954 => x"3367d700",
         955 => x"93060e00",
         956 => x"637e0701",
         957 => x"3307e500",
         958 => x"9306feff",
         959 => x"6368a700",
         960 => x"63760701",
         961 => x"9306eeff",
         962 => x"3307a700",
         963 => x"93970701",
         964 => x"33e5d700",
         965 => x"13130601",
         966 => x"93960601",
         967 => x"93d60601",
         968 => x"13530301",
         969 => x"13560601",
         970 => x"33070741",
         971 => x"13580501",
         972 => x"338e6602",
         973 => x"33036802",
         974 => x"93570e01",
         975 => x"b386c602",
         976 => x"b3866600",
         977 => x"b387d700",
         978 => x"3308c802",
         979 => x"63f66700",
         980 => x"b7060100",
         981 => x"3308d800",
         982 => x"93d60701",
         983 => x"b3860601",
         984 => x"6362d702",
         985 => x"e31cd7ce",
         986 => x"131e0e01",
         987 => x"93970701",
         988 => x"135e0e01",
         989 => x"b398b800",
         990 => x"b387c701",
         991 => x"93050000",
         992 => x"e3f0f8ce",
         993 => x"1305f5ff",
         994 => x"6ff05fcd",
         995 => x"93050000",
         996 => x"13050000",
         997 => x"67800000",
         998 => x"13080600",
         999 => x"93070500",
        1000 => x"13870500",
        1001 => x"63960620",
        1002 => x"b7380000",
        1003 => x"9388c8b6",
        1004 => x"63fcc50c",
        1005 => x"b7060100",
        1006 => x"637ed60a",
        1007 => x"93360610",
        1008 => x"93b61600",
        1009 => x"93963600",
        1010 => x"3353d600",
        1011 => x"b3886800",
        1012 => x"83c80800",
        1013 => x"13030002",
        1014 => x"b386d800",
        1015 => x"b308d340",
        1016 => x"630cd300",
        1017 => x"33971501",
        1018 => x"b356d500",
        1019 => x"33181601",
        1020 => x"33e7e600",
        1021 => x"b3171501",
        1022 => x"13560801",
        1023 => x"b356c702",
        1024 => x"13150801",
        1025 => x"13550501",
        1026 => x"3377c702",
        1027 => x"b386a602",
        1028 => x"93150701",
        1029 => x"13d70701",
        1030 => x"3367b700",
        1031 => x"637ad700",
        1032 => x"3307e800",
        1033 => x"63660701",
        1034 => x"6374d700",
        1035 => x"33070701",
        1036 => x"3307d740",
        1037 => x"b356c702",
        1038 => x"3377c702",
        1039 => x"b386a602",
        1040 => x"93970701",
        1041 => x"13170701",
        1042 => x"93d70701",
        1043 => x"b3e7e700",
        1044 => x"63fad700",
        1045 => x"b307f800",
        1046 => x"63e60701",
        1047 => x"63f4d700",
        1048 => x"b3870701",
        1049 => x"b387d740",
        1050 => x"33d51701",
        1051 => x"93050000",
        1052 => x"67800000",
        1053 => x"37030001",
        1054 => x"93068001",
        1055 => x"e37666f4",
        1056 => x"93060001",
        1057 => x"6ff05ff4",
        1058 => x"93060000",
        1059 => x"630c0600",
        1060 => x"37070100",
        1061 => x"637ee606",
        1062 => x"93360610",
        1063 => x"93b61600",
        1064 => x"93963600",
        1065 => x"3357d600",
        1066 => x"b388e800",
        1067 => x"03c70800",
        1068 => x"3307d700",
        1069 => x"93060002",
        1070 => x"b388e640",
        1071 => x"6394e606",
        1072 => x"3387c540",
        1073 => x"93550801",
        1074 => x"3356b702",
        1075 => x"13150801",
        1076 => x"13550501",
        1077 => x"93d60701",
        1078 => x"3377b702",
        1079 => x"3306a602",
        1080 => x"13170701",
        1081 => x"33e7e600",
        1082 => x"637ac700",
        1083 => x"3307e800",
        1084 => x"63660701",
        1085 => x"6374c700",
        1086 => x"33070701",
        1087 => x"3307c740",
        1088 => x"b356b702",
        1089 => x"3377b702",
        1090 => x"b386a602",
        1091 => x"6ff05ff3",
        1092 => x"37070001",
        1093 => x"93068001",
        1094 => x"e376e6f8",
        1095 => x"93060001",
        1096 => x"6ff05ff8",
        1097 => x"33181601",
        1098 => x"b3d6e500",
        1099 => x"b3171501",
        1100 => x"b3951501",
        1101 => x"3357e500",
        1102 => x"13550801",
        1103 => x"3367b700",
        1104 => x"b3d5a602",
        1105 => x"13130801",
        1106 => x"13530301",
        1107 => x"b3f6a602",
        1108 => x"b3856502",
        1109 => x"13960601",
        1110 => x"93560701",
        1111 => x"b3e6c600",
        1112 => x"63fab600",
        1113 => x"b306d800",
        1114 => x"63e60601",
        1115 => x"63f4b600",
        1116 => x"b3860601",
        1117 => x"b386b640",
        1118 => x"33d6a602",
        1119 => x"13170701",
        1120 => x"13570701",
        1121 => x"b3f6a602",
        1122 => x"33066602",
        1123 => x"93960601",
        1124 => x"3367d700",
        1125 => x"637ac700",
        1126 => x"3307e800",
        1127 => x"63660701",
        1128 => x"6374c700",
        1129 => x"33070701",
        1130 => x"3307c740",
        1131 => x"6ff09ff1",
        1132 => x"63e2d51c",
        1133 => x"37080100",
        1134 => x"63fe0605",
        1135 => x"13b80610",
        1136 => x"13381800",
        1137 => x"13183800",
        1138 => x"b7380000",
        1139 => x"33d30601",
        1140 => x"9388c8b6",
        1141 => x"b3886800",
        1142 => x"83c80800",
        1143 => x"13030002",
        1144 => x"b3880801",
        1145 => x"33081341",
        1146 => x"63101305",
        1147 => x"63e4b600",
        1148 => x"636cc500",
        1149 => x"3306c540",
        1150 => x"b386d540",
        1151 => x"3337c500",
        1152 => x"93070600",
        1153 => x"3387e640",
        1154 => x"13850700",
        1155 => x"93050700",
        1156 => x"67800000",
        1157 => x"b7080001",
        1158 => x"13088001",
        1159 => x"e3f616fb",
        1160 => x"13080001",
        1161 => x"6ff05ffa",
        1162 => x"b3571601",
        1163 => x"b3960601",
        1164 => x"b3e6d700",
        1165 => x"33d71501",
        1166 => x"13d30601",
        1167 => x"335f6702",
        1168 => x"139e0601",
        1169 => x"135e0e01",
        1170 => x"b3970501",
        1171 => x"b3551501",
        1172 => x"b3e5f500",
        1173 => x"93d70501",
        1174 => x"33160601",
        1175 => x"33150501",
        1176 => x"33776702",
        1177 => x"b30eee03",
        1178 => x"13170701",
        1179 => x"b3e7e700",
        1180 => x"13070f00",
        1181 => x"63fed701",
        1182 => x"b387f600",
        1183 => x"1307ffff",
        1184 => x"63e8d700",
        1185 => x"63f6d701",
        1186 => x"1307efff",
        1187 => x"b387d700",
        1188 => x"b387d741",
        1189 => x"b3de6702",
        1190 => x"93950501",
        1191 => x"93d50501",
        1192 => x"b3f76702",
        1193 => x"13830e00",
        1194 => x"330ede03",
        1195 => x"93970701",
        1196 => x"b3e5f500",
        1197 => x"63fec501",
        1198 => x"b385b600",
        1199 => x"1383feff",
        1200 => x"63e8d500",
        1201 => x"63f6c501",
        1202 => x"1383eeff",
        1203 => x"b385d500",
        1204 => x"93170701",
        1205 => x"b3e76700",
        1206 => x"b385c541",
        1207 => x"13130301",
        1208 => x"131e0601",
        1209 => x"13570601",
        1210 => x"13530301",
        1211 => x"93d70701",
        1212 => x"135e0e01",
        1213 => x"b30ec303",
        1214 => x"338ec703",
        1215 => x"3303e302",
        1216 => x"b387e702",
        1217 => x"3303c301",
        1218 => x"13d70e01",
        1219 => x"33076700",
        1220 => x"6376c701",
        1221 => x"37030100",
        1222 => x"b3876700",
        1223 => x"13530701",
        1224 => x"939e0e01",
        1225 => x"13170701",
        1226 => x"93de0e01",
        1227 => x"b307f300",
        1228 => x"3307d701",
        1229 => x"63e6f500",
        1230 => x"639ef500",
        1231 => x"637ce500",
        1232 => x"3306c740",
        1233 => x"3333c700",
        1234 => x"b306d300",
        1235 => x"13070600",
        1236 => x"b387d740",
        1237 => x"3307e540",
        1238 => x"3335e500",
        1239 => x"b385f540",
        1240 => x"b385a540",
        1241 => x"b3981501",
        1242 => x"33570701",
        1243 => x"33e5e800",
        1244 => x"b3d50501",
        1245 => x"67800000",
        1246 => x"13030500",
        1247 => x"630a0600",
        1248 => x"2300b300",
        1249 => x"1306f6ff",
        1250 => x"13031300",
        1251 => x"e31a06fe",
        1252 => x"67800000",
        1253 => x"13030500",
        1254 => x"630e0600",
        1255 => x"83830500",
        1256 => x"23007300",
        1257 => x"1306f6ff",
        1258 => x"13031300",
        1259 => x"93851500",
        1260 => x"e31606fe",
        1261 => x"67800000",
        1262 => x"630c0602",
        1263 => x"13030500",
        1264 => x"93061000",
        1265 => x"636ab500",
        1266 => x"9306f0ff",
        1267 => x"1307f6ff",
        1268 => x"3303e300",
        1269 => x"b385e500",
        1270 => x"83830500",
        1271 => x"23007300",
        1272 => x"1306f6ff",
        1273 => x"3303d300",
        1274 => x"b385d500",
        1275 => x"e31606fe",
        1276 => x"67800000",
        1277 => x"6f000000",
        1278 => x"130101ff",
        1279 => x"23248100",
        1280 => x"13040000",
        1281 => x"23229100",
        1282 => x"23202101",
        1283 => x"23261100",
        1284 => x"93040500",
        1285 => x"13090400",
        1286 => x"93070400",
        1287 => x"732410c8",
        1288 => x"732910c0",
        1289 => x"f32710c8",
        1290 => x"e31af4fe",
        1291 => x"37460f00",
        1292 => x"13060624",
        1293 => x"93060000",
        1294 => x"13050900",
        1295 => x"93050400",
        1296 => x"eff09fb5",
        1297 => x"37460f00",
        1298 => x"23a4a400",
        1299 => x"93050400",
        1300 => x"13050900",
        1301 => x"13060624",
        1302 => x"93060000",
        1303 => x"eff00ff1",
        1304 => x"8320c100",
        1305 => x"03248100",
        1306 => x"23a0a400",
        1307 => x"23a2b400",
        1308 => x"03290100",
        1309 => x"83244100",
        1310 => x"13050000",
        1311 => x"13010101",
        1312 => x"67800000",
        1313 => x"03a78186",
        1314 => x"b7870020",
        1315 => x"93870700",
        1316 => x"93060040",
        1317 => x"b387d740",
        1318 => x"630c0700",
        1319 => x"3305a700",
        1320 => x"63e2a702",
        1321 => x"23a4a186",
        1322 => x"13050700",
        1323 => x"67800000",
        1324 => x"9386819b",
        1325 => x"1387819b",
        1326 => x"23a4d186",
        1327 => x"3305a700",
        1328 => x"e3f2a7fe",
        1329 => x"130101ff",
        1330 => x"23261100",
        1331 => x"ef00c054",
        1332 => x"8320c100",
        1333 => x"9307c000",
        1334 => x"2320f500",
        1335 => x"1307f0ff",
        1336 => x"13050700",
        1337 => x"13010101",
        1338 => x"67800000",
        1339 => x"370700f0",
        1340 => x"13070710",
        1341 => x"83274700",
        1342 => x"93f78700",
        1343 => x"e38c07fe",
        1344 => x"03258700",
        1345 => x"1375f50f",
        1346 => x"67800000",
        1347 => x"f32710fc",
        1348 => x"63960700",
        1349 => x"b7f7fa02",
        1350 => x"93870708",
        1351 => x"63060500",
        1352 => x"33d5a702",
        1353 => x"1305f5ff",
        1354 => x"b70700f0",
        1355 => x"23a6a710",
        1356 => x"23a0b710",
        1357 => x"23a20710",
        1358 => x"67800000",
        1359 => x"370700f0",
        1360 => x"1375f50f",
        1361 => x"13070710",
        1362 => x"2324a700",
        1363 => x"83274700",
        1364 => x"93f70701",
        1365 => x"e38c07fe",
        1366 => x"67800000",
        1367 => x"630e0502",
        1368 => x"130101ff",
        1369 => x"23248100",
        1370 => x"23261100",
        1371 => x"13040500",
        1372 => x"03450500",
        1373 => x"630a0500",
        1374 => x"13041400",
        1375 => x"eff01ffc",
        1376 => x"03450400",
        1377 => x"e31a05fe",
        1378 => x"8320c100",
        1379 => x"03248100",
        1380 => x"13010101",
        1381 => x"67800000",
        1382 => x"67800000",
        1383 => x"130101f9",
        1384 => x"23229106",
        1385 => x"23202107",
        1386 => x"23261106",
        1387 => x"23248106",
        1388 => x"232e3105",
        1389 => x"232c4105",
        1390 => x"232a5105",
        1391 => x"23286105",
        1392 => x"23267105",
        1393 => x"23248105",
        1394 => x"23229105",
        1395 => x"13090500",
        1396 => x"93840500",
        1397 => x"f32a00fc",
        1398 => x"b7070008",
        1399 => x"232c0100",
        1400 => x"232e0100",
        1401 => x"23200102",
        1402 => x"23220102",
        1403 => x"23240102",
        1404 => x"23260102",
        1405 => x"23280102",
        1406 => x"232a0102",
        1407 => x"232c0102",
        1408 => x"232e0102",
        1409 => x"b3fafa00",
        1410 => x"732410fc",
        1411 => x"63160400",
        1412 => x"37f4fa02",
        1413 => x"13040408",
        1414 => x"97f2ffff",
        1415 => x"938282ce",
        1416 => x"73905230",
        1417 => x"37c50100",
        1418 => x"13050520",
        1419 => x"93059000",
        1420 => x"eff0dfed",
        1421 => x"b717b7d1",
        1422 => x"93879775",
        1423 => x"b337f402",
        1424 => x"93561400",
        1425 => x"37353e05",
        1426 => x"370600f0",
        1427 => x"13576400",
        1428 => x"130535d6",
        1429 => x"9386f6ff",
        1430 => x"2326d660",
        1431 => x"b725d96f",
        1432 => x"93060600",
        1433 => x"3337a702",
        1434 => x"93d7d700",
        1435 => x"13051001",
        1436 => x"2320a660",
        1437 => x"938555d8",
        1438 => x"9387f7ff",
        1439 => x"23a8f670",
        1440 => x"37260000",
        1441 => x"1306f670",
        1442 => x"23a6c670",
        1443 => x"b337b402",
        1444 => x"13576700",
        1445 => x"1307f7ff",
        1446 => x"23a0a670",
        1447 => x"93058070",
        1448 => x"13170701",
        1449 => x"23a0b640",
        1450 => x"13678700",
        1451 => x"23a0e620",
        1452 => x"1307a007",
        1453 => x"93d73701",
        1454 => x"9387f7ff",
        1455 => x"93970701",
        1456 => x"93e7c700",
        1457 => x"23a0f630",
        1458 => x"23ace600",
        1459 => x"f3224030",
        1460 => x"93e20208",
        1461 => x"73904230",
        1462 => x"f3224030",
        1463 => x"93e28200",
        1464 => x"73904230",
        1465 => x"b7220000",
        1466 => x"93828280",
        1467 => x"73900230",
        1468 => x"b7390000",
        1469 => x"1385c9c8",
        1470 => x"eff05fe6",
        1471 => x"1304f9ff",
        1472 => x"63522003",
        1473 => x"1309f0ff",
        1474 => x"03a50400",
        1475 => x"1304f4ff",
        1476 => x"93844400",
        1477 => x"eff09fe4",
        1478 => x"1385c9c8",
        1479 => x"eff01fe4",
        1480 => x"e31424ff",
        1481 => x"37350000",
        1482 => x"130505c9",
        1483 => x"eff01fe3",
        1484 => x"63960a22",
        1485 => x"b7040010",
        1486 => x"b7998888",
        1487 => x"37f4eeee",
        1488 => x"9384f4ff",
        1489 => x"93899988",
        1490 => x"1304f4ee",
        1491 => x"373a0000",
        1492 => x"b71b0000",
        1493 => x"37f9eeee",
        1494 => x"938b0b2c",
        1495 => x"1309e9ee",
        1496 => x"6f00c000",
        1497 => x"938bfbff",
        1498 => x"63860b1a",
        1499 => x"93050000",
        1500 => x"13058100",
        1501 => x"ef008034",
        1502 => x"e31605fe",
        1503 => x"032c8100",
        1504 => x"8325c100",
        1505 => x"37160000",
        1506 => x"9357cc01",
        1507 => x"13974500",
        1508 => x"b367f700",
        1509 => x"33f79700",
        1510 => x"b3779c00",
        1511 => x"13d58501",
        1512 => x"b387e700",
        1513 => x"13d7f541",
        1514 => x"b387a700",
        1515 => x"1375d700",
        1516 => x"b387a700",
        1517 => x"33b83703",
        1518 => x"137727ff",
        1519 => x"130606e1",
        1520 => x"93060000",
        1521 => x"13050c00",
        1522 => x"938bfbff",
        1523 => x"13583800",
        1524 => x"93184800",
        1525 => x"33880841",
        1526 => x"b3870741",
        1527 => x"b387e700",
        1528 => x"13d7f741",
        1529 => x"b307fc40",
        1530 => x"3338fc00",
        1531 => x"3387e540",
        1532 => x"33070741",
        1533 => x"b3882703",
        1534 => x"33078702",
        1535 => x"33b88702",
        1536 => x"33071701",
        1537 => x"b3878702",
        1538 => x"33070701",
        1539 => x"1358f741",
        1540 => x"13783800",
        1541 => x"b307f800",
        1542 => x"33b80701",
        1543 => x"3308e800",
        1544 => x"1317e801",
        1545 => x"93d72700",
        1546 => x"b367f700",
        1547 => x"93582840",
        1548 => x"13d7c701",
        1549 => x"13934800",
        1550 => x"3367e300",
        1551 => x"33739700",
        1552 => x"33f79700",
        1553 => x"1358f841",
        1554 => x"33076700",
        1555 => x"13d38801",
        1556 => x"33076700",
        1557 => x"1373d800",
        1558 => x"33076700",
        1559 => x"33333703",
        1560 => x"137828ff",
        1561 => x"139b4700",
        1562 => x"330bfb40",
        1563 => x"131b2b00",
        1564 => x"330b6c41",
        1565 => x"13533300",
        1566 => x"131e4300",
        1567 => x"33036e40",
        1568 => x"33076740",
        1569 => x"33070701",
        1570 => x"1358f741",
        1571 => x"3387e740",
        1572 => x"33880841",
        1573 => x"b3b8e700",
        1574 => x"33081841",
        1575 => x"33032703",
        1576 => x"33088802",
        1577 => x"b3388702",
        1578 => x"33086800",
        1579 => x"33078702",
        1580 => x"33081801",
        1581 => x"9358f841",
        1582 => x"93f83800",
        1583 => x"3387e800",
        1584 => x"b3381701",
        1585 => x"b3880801",
        1586 => x"9398e801",
        1587 => x"13572700",
        1588 => x"33e7e800",
        1589 => x"13184700",
        1590 => x"3307e840",
        1591 => x"13172700",
        1592 => x"b38ce740",
        1593 => x"efe05fe1",
        1594 => x"83260101",
        1595 => x"13070500",
        1596 => x"13080b00",
        1597 => x"93870c00",
        1598 => x"13060c00",
        1599 => x"93058acf",
        1600 => x"13058101",
        1601 => x"ef00000a",
        1602 => x"13058101",
        1603 => x"eff01fc5",
        1604 => x"e39e0be4",
        1605 => x"63940a00",
        1606 => x"73001000",
        1607 => x"b70700f0",
        1608 => x"9306f00f",
        1609 => x"23a4d740",
        1610 => x"83a60720",
        1611 => x"13060009",
        1612 => x"371700f0",
        1613 => x"93e60630",
        1614 => x"23a0d720",
        1615 => x"23a4c720",
        1616 => x"83a60730",
        1617 => x"93e60630",
        1618 => x"23a0d730",
        1619 => x"23a4c730",
        1620 => x"93071000",
        1621 => x"2320f790",
        1622 => x"6ff09fdf",
        1623 => x"37350000",
        1624 => x"130505cc",
        1625 => x"eff09fbf",
        1626 => x"6ff0dfdc",
        1627 => x"130101ff",
        1628 => x"23248100",
        1629 => x"23261100",
        1630 => x"93070000",
        1631 => x"13040500",
        1632 => x"63880700",
        1633 => x"93050000",
        1634 => x"97000000",
        1635 => x"e7000000",
        1636 => x"83a7c186",
        1637 => x"63840700",
        1638 => x"e7800700",
        1639 => x"13050400",
        1640 => x"eff05fa5",
        1641 => x"130101f6",
        1642 => x"232af108",
        1643 => x"b7070080",
        1644 => x"9387f7ff",
        1645 => x"232ef100",
        1646 => x"2328f100",
        1647 => x"b707ffff",
        1648 => x"93878720",
        1649 => x"232af100",
        1650 => x"2324a100",
        1651 => x"232ca100",
        1652 => x"03a54186",
        1653 => x"2324c108",
        1654 => x"2326d108",
        1655 => x"13860500",
        1656 => x"93068108",
        1657 => x"93058100",
        1658 => x"232e1106",
        1659 => x"2328e108",
        1660 => x"232c0109",
        1661 => x"232e1109",
        1662 => x"23260106",
        1663 => x"2322d100",
        1664 => x"ef000058",
        1665 => x"83278100",
        1666 => x"23800700",
        1667 => x"8320c107",
        1668 => x"1301010a",
        1669 => x"67800000",
        1670 => x"03a54186",
        1671 => x"67800000",
        1672 => x"130101ff",
        1673 => x"23248100",
        1674 => x"23229100",
        1675 => x"37340000",
        1676 => x"b7340000",
        1677 => x"938784e5",
        1678 => x"130484e5",
        1679 => x"3304f440",
        1680 => x"23202101",
        1681 => x"23261100",
        1682 => x"13542440",
        1683 => x"938484e5",
        1684 => x"13090000",
        1685 => x"63108904",
        1686 => x"b7340000",
        1687 => x"37340000",
        1688 => x"938784e5",
        1689 => x"130484e5",
        1690 => x"3304f440",
        1691 => x"13542440",
        1692 => x"938484e5",
        1693 => x"13090000",
        1694 => x"63188902",
        1695 => x"8320c100",
        1696 => x"03248100",
        1697 => x"83244100",
        1698 => x"03290100",
        1699 => x"13010101",
        1700 => x"67800000",
        1701 => x"83a70400",
        1702 => x"13091900",
        1703 => x"93844400",
        1704 => x"e7800700",
        1705 => x"6ff01ffb",
        1706 => x"83a70400",
        1707 => x"13091900",
        1708 => x"93844400",
        1709 => x"e7800700",
        1710 => x"6ff01ffc",
        1711 => x"13860500",
        1712 => x"93050500",
        1713 => x"03a54186",
        1714 => x"6f00105a",
        1715 => x"638a050e",
        1716 => x"83a7c5ff",
        1717 => x"130101fe",
        1718 => x"232c8100",
        1719 => x"232e1100",
        1720 => x"1384c5ff",
        1721 => x"63d40700",
        1722 => x"3304f400",
        1723 => x"2326a100",
        1724 => x"ef004031",
        1725 => x"83a78187",
        1726 => x"0325c100",
        1727 => x"639e0700",
        1728 => x"23220400",
        1729 => x"23ac8186",
        1730 => x"03248101",
        1731 => x"8320c101",
        1732 => x"13010102",
        1733 => x"6f00402f",
        1734 => x"6374f402",
        1735 => x"03260400",
        1736 => x"b306c400",
        1737 => x"639ad700",
        1738 => x"83a60700",
        1739 => x"83a74700",
        1740 => x"b386c600",
        1741 => x"2320d400",
        1742 => x"2322f400",
        1743 => x"6ff09ffc",
        1744 => x"13870700",
        1745 => x"83a74700",
        1746 => x"63840700",
        1747 => x"e37af4fe",
        1748 => x"83260700",
        1749 => x"3306d700",
        1750 => x"63188602",
        1751 => x"03260400",
        1752 => x"b386c600",
        1753 => x"2320d700",
        1754 => x"3306d700",
        1755 => x"e39ec7f8",
        1756 => x"03a60700",
        1757 => x"83a74700",
        1758 => x"b306d600",
        1759 => x"2320d700",
        1760 => x"2322f700",
        1761 => x"6ff05ff8",
        1762 => x"6378c400",
        1763 => x"9307c000",
        1764 => x"2320f500",
        1765 => x"6ff05ff7",
        1766 => x"03260400",
        1767 => x"b306c400",
        1768 => x"639ad700",
        1769 => x"83a60700",
        1770 => x"83a74700",
        1771 => x"b386c600",
        1772 => x"2320d400",
        1773 => x"2322f400",
        1774 => x"23228700",
        1775 => x"6ff0dff4",
        1776 => x"67800000",
        1777 => x"130101ff",
        1778 => x"23202101",
        1779 => x"83a74187",
        1780 => x"23248100",
        1781 => x"23229100",
        1782 => x"23261100",
        1783 => x"93040500",
        1784 => x"13840500",
        1785 => x"63980700",
        1786 => x"93050000",
        1787 => x"ef00904c",
        1788 => x"23aaa186",
        1789 => x"93050400",
        1790 => x"13850400",
        1791 => x"ef00904b",
        1792 => x"1309f0ff",
        1793 => x"63122503",
        1794 => x"1304f0ff",
        1795 => x"8320c100",
        1796 => x"13050400",
        1797 => x"03248100",
        1798 => x"83244100",
        1799 => x"03290100",
        1800 => x"13010101",
        1801 => x"67800000",
        1802 => x"13043500",
        1803 => x"1374c4ff",
        1804 => x"e30e85fc",
        1805 => x"b305a440",
        1806 => x"13850400",
        1807 => x"ef009047",
        1808 => x"e31625fd",
        1809 => x"6ff05ffc",
        1810 => x"130101fe",
        1811 => x"232a9100",
        1812 => x"93843500",
        1813 => x"93f4c4ff",
        1814 => x"23282101",
        1815 => x"232e1100",
        1816 => x"232c8100",
        1817 => x"23263101",
        1818 => x"23244101",
        1819 => x"93848400",
        1820 => x"9307c000",
        1821 => x"13090500",
        1822 => x"63fef408",
        1823 => x"93840700",
        1824 => x"63ecb408",
        1825 => x"13050900",
        1826 => x"ef00c017",
        1827 => x"83a78187",
        1828 => x"13840700",
        1829 => x"6316040a",
        1830 => x"93850400",
        1831 => x"13050900",
        1832 => x"eff05ff2",
        1833 => x"9307f0ff",
        1834 => x"13040500",
        1835 => x"6318f514",
        1836 => x"03a48187",
        1837 => x"93070400",
        1838 => x"63980710",
        1839 => x"63060412",
        1840 => x"032a0400",
        1841 => x"93050000",
        1842 => x"13050900",
        1843 => x"330a4401",
        1844 => x"ef00503e",
        1845 => x"631aaa10",
        1846 => x"83270400",
        1847 => x"13050900",
        1848 => x"b384f440",
        1849 => x"93850400",
        1850 => x"eff0dfed",
        1851 => x"9307f0ff",
        1852 => x"630cf50e",
        1853 => x"83270400",
        1854 => x"b3879700",
        1855 => x"2320f400",
        1856 => x"83a78187",
        1857 => x"03a74700",
        1858 => x"6316070c",
        1859 => x"23ac0186",
        1860 => x"6f000006",
        1861 => x"e3d604f6",
        1862 => x"2320f900",
        1863 => x"13050000",
        1864 => x"8320c101",
        1865 => x"03248101",
        1866 => x"83244101",
        1867 => x"03290101",
        1868 => x"8329c100",
        1869 => x"032a8100",
        1870 => x"13010102",
        1871 => x"67800000",
        1872 => x"83260400",
        1873 => x"b3869640",
        1874 => x"63ca0606",
        1875 => x"1307b000",
        1876 => x"637ad704",
        1877 => x"23209400",
        1878 => x"33079400",
        1879 => x"63908704",
        1880 => x"23ace186",
        1881 => x"83274400",
        1882 => x"2320d700",
        1883 => x"2322f700",
        1884 => x"13050900",
        1885 => x"ef004009",
        1886 => x"1305b400",
        1887 => x"93074400",
        1888 => x"137585ff",
        1889 => x"3307f540",
        1890 => x"e30cf5f8",
        1891 => x"3304e400",
        1892 => x"b387a740",
        1893 => x"2320f400",
        1894 => x"6ff09ff8",
        1895 => x"23a2e700",
        1896 => x"6ff05ffc",
        1897 => x"03274400",
        1898 => x"63968700",
        1899 => x"23ace186",
        1900 => x"6ff01ffc",
        1901 => x"23a2e700",
        1902 => x"6ff09ffb",
        1903 => x"93070400",
        1904 => x"03244400",
        1905 => x"6ff01fed",
        1906 => x"13840700",
        1907 => x"83a74700",
        1908 => x"6ff09fee",
        1909 => x"13870700",
        1910 => x"83a74700",
        1911 => x"e39c87fe",
        1912 => x"23220700",
        1913 => x"6ff0dff8",
        1914 => x"9307c000",
        1915 => x"2320f900",
        1916 => x"13050900",
        1917 => x"ef004001",
        1918 => x"6ff05ff2",
        1919 => x"23209500",
        1920 => x"6ff01ff7",
        1921 => x"67800000",
        1922 => x"67800000",
        1923 => x"130101fe",
        1924 => x"23282101",
        1925 => x"03a98500",
        1926 => x"232c8100",
        1927 => x"23263101",
        1928 => x"23244101",
        1929 => x"232e1100",
        1930 => x"232a9100",
        1931 => x"23225101",
        1932 => x"23206101",
        1933 => x"13840500",
        1934 => x"130a0600",
        1935 => x"93890600",
        1936 => x"63ec2613",
        1937 => x"8397c500",
        1938 => x"13070900",
        1939 => x"93f60748",
        1940 => x"638c0608",
        1941 => x"83244401",
        1942 => x"13073000",
        1943 => x"83a50501",
        1944 => x"b384e402",
        1945 => x"13072000",
        1946 => x"832a0400",
        1947 => x"130b0500",
        1948 => x"b38aba40",
        1949 => x"b3c4e402",
        1950 => x"13871900",
        1951 => x"33075701",
        1952 => x"13860400",
        1953 => x"63f6e400",
        1954 => x"93040700",
        1955 => x"13060700",
        1956 => x"93f70740",
        1957 => x"6386070a",
        1958 => x"93050600",
        1959 => x"13050b00",
        1960 => x"eff09fda",
        1961 => x"13090500",
        1962 => x"630a050a",
        1963 => x"83250401",
        1964 => x"13860a00",
        1965 => x"eff00fce",
        1966 => x"8357c400",
        1967 => x"93f7f7b7",
        1968 => x"93e70708",
        1969 => x"2316f400",
        1970 => x"23282401",
        1971 => x"232a9400",
        1972 => x"33095901",
        1973 => x"b3845441",
        1974 => x"23202401",
        1975 => x"23249400",
        1976 => x"13890900",
        1977 => x"13870900",
        1978 => x"93090700",
        1979 => x"03250400",
        1980 => x"13860900",
        1981 => x"93050a00",
        1982 => x"eff00fcc",
        1983 => x"83278400",
        1984 => x"13050000",
        1985 => x"b3872741",
        1986 => x"2324f400",
        1987 => x"83270400",
        1988 => x"b3873701",
        1989 => x"2320f400",
        1990 => x"8320c101",
        1991 => x"03248101",
        1992 => x"83244101",
        1993 => x"03290101",
        1994 => x"8329c100",
        1995 => x"032a8100",
        1996 => x"832a4100",
        1997 => x"032b0100",
        1998 => x"13010102",
        1999 => x"67800000",
        2000 => x"13050b00",
        2001 => x"ef00901b",
        2002 => x"13090500",
        2003 => x"e31e05f6",
        2004 => x"83250401",
        2005 => x"13050b00",
        2006 => x"eff05fb7",
        2007 => x"9307c000",
        2008 => x"2320fb00",
        2009 => x"8357c400",
        2010 => x"1305f0ff",
        2011 => x"93e70704",
        2012 => x"2316f400",
        2013 => x"6ff05ffa",
        2014 => x"13890600",
        2015 => x"6ff01ff7",
        2016 => x"83d7c500",
        2017 => x"130101f6",
        2018 => x"232c8108",
        2019 => x"232a9108",
        2020 => x"23282109",
        2021 => x"23244109",
        2022 => x"232e1108",
        2023 => x"23263109",
        2024 => x"23225109",
        2025 => x"23206109",
        2026 => x"232e7107",
        2027 => x"232c8107",
        2028 => x"232a9107",
        2029 => x"93f70708",
        2030 => x"130a0500",
        2031 => x"13890500",
        2032 => x"93040600",
        2033 => x"13840600",
        2034 => x"63840706",
        2035 => x"83a70501",
        2036 => x"63900706",
        2037 => x"93050004",
        2038 => x"eff01fc7",
        2039 => x"2320a900",
        2040 => x"2328a900",
        2041 => x"63120504",
        2042 => x"9307c000",
        2043 => x"2320fa00",
        2044 => x"1305f0ff",
        2045 => x"8320c109",
        2046 => x"03248109",
        2047 => x"83244109",
        2048 => x"03290109",
        2049 => x"8329c108",
        2050 => x"032a8108",
        2051 => x"832a4108",
        2052 => x"032b0108",
        2053 => x"832bc107",
        2054 => x"032c8107",
        2055 => x"832c4107",
        2056 => x"1301010a",
        2057 => x"67800000",
        2058 => x"93070004",
        2059 => x"232af900",
        2060 => x"93070002",
        2061 => x"a304f102",
        2062 => x"93070003",
        2063 => x"23220102",
        2064 => x"2305f102",
        2065 => x"23268100",
        2066 => x"930b5002",
        2067 => x"930af0ff",
        2068 => x"130c1000",
        2069 => x"130ba000",
        2070 => x"13840400",
        2071 => x"83470400",
        2072 => x"63840700",
        2073 => x"6396770d",
        2074 => x"b30c9440",
        2075 => x"63049402",
        2076 => x"93860c00",
        2077 => x"13860400",
        2078 => x"93050900",
        2079 => x"13050a00",
        2080 => x"eff0dfd8",
        2081 => x"63045525",
        2082 => x"83274102",
        2083 => x"b3879701",
        2084 => x"2322f102",
        2085 => x"83470400",
        2086 => x"638a0722",
        2087 => x"93041400",
        2088 => x"23280100",
        2089 => x"232e0100",
        2090 => x"232a5101",
        2091 => x"232c0100",
        2092 => x"a3090104",
        2093 => x"23240106",
        2094 => x"b73c0000",
        2095 => x"83c50400",
        2096 => x"13065000",
        2097 => x"13854cdc",
        2098 => x"ef00c077",
        2099 => x"03270101",
        2100 => x"93070500",
        2101 => x"13841400",
        2102 => x"63100506",
        2103 => x"93770701",
        2104 => x"63860700",
        2105 => x"93070002",
        2106 => x"a309f104",
        2107 => x"93778700",
        2108 => x"63860700",
        2109 => x"9307b002",
        2110 => x"a309f104",
        2111 => x"83c60400",
        2112 => x"9307a002",
        2113 => x"6388f604",
        2114 => x"8327c101",
        2115 => x"13840400",
        2116 => x"93060000",
        2117 => x"13069000",
        2118 => x"03470400",
        2119 => x"93051400",
        2120 => x"130707fd",
        2121 => x"637ce608",
        2122 => x"63900604",
        2123 => x"6f004005",
        2124 => x"13041400",
        2125 => x"6ff09ff2",
        2126 => x"93864cdc",
        2127 => x"b387d740",
        2128 => x"b317fc00",
        2129 => x"b3e7e700",
        2130 => x"2328f100",
        2131 => x"93040400",
        2132 => x"6ff0dff6",
        2133 => x"8327c100",
        2134 => x"93864700",
        2135 => x"83a70700",
        2136 => x"2326d100",
        2137 => x"63c60700",
        2138 => x"232ef100",
        2139 => x"6f004001",
        2140 => x"b307f040",
        2141 => x"13672700",
        2142 => x"232ef100",
        2143 => x"2328e100",
        2144 => x"03470400",
        2145 => x"9307e002",
        2146 => x"6318f706",
        2147 => x"03471400",
        2148 => x"9307a002",
        2149 => x"631ef702",
        2150 => x"8327c100",
        2151 => x"13042400",
        2152 => x"13874700",
        2153 => x"83a70700",
        2154 => x"2326e100",
        2155 => x"63d40700",
        2156 => x"9307f0ff",
        2157 => x"232af100",
        2158 => x"6f000004",
        2159 => x"b3876703",
        2160 => x"13840500",
        2161 => x"93061000",
        2162 => x"b387e700",
        2163 => x"6ff0dff4",
        2164 => x"13041400",
        2165 => x"232a0100",
        2166 => x"93060000",
        2167 => x"93070000",
        2168 => x"13069000",
        2169 => x"03470400",
        2170 => x"93051400",
        2171 => x"130707fd",
        2172 => x"6378e608",
        2173 => x"e39006fc",
        2174 => x"83450400",
        2175 => x"b7340000",
        2176 => x"13063000",
        2177 => x"1385c4dc",
        2178 => x"ef00c063",
        2179 => x"63020502",
        2180 => x"83270101",
        2181 => x"9384c4dc",
        2182 => x"33059540",
        2183 => x"13070004",
        2184 => x"3317a700",
        2185 => x"b3e7e700",
        2186 => x"13041400",
        2187 => x"2328f100",
        2188 => x"83450400",
        2189 => x"37350000",
        2190 => x"13066000",
        2191 => x"130505dd",
        2192 => x"93041400",
        2193 => x"2304b102",
        2194 => x"ef00c05f",
        2195 => x"630a0508",
        2196 => x"93070000",
        2197 => x"63980704",
        2198 => x"03270101",
        2199 => x"8327c100",
        2200 => x"13770710",
        2201 => x"63080702",
        2202 => x"93874700",
        2203 => x"2326f100",
        2204 => x"83274102",
        2205 => x"b3873701",
        2206 => x"2322f102",
        2207 => x"6ff0dfdd",
        2208 => x"b3876703",
        2209 => x"13840500",
        2210 => x"93061000",
        2211 => x"b387e700",
        2212 => x"6ff05ff5",
        2213 => x"93877700",
        2214 => x"93f787ff",
        2215 => x"93878700",
        2216 => x"6ff0dffc",
        2217 => x"b7260000",
        2218 => x"1307c100",
        2219 => x"9386c6e0",
        2220 => x"13060900",
        2221 => x"93050101",
        2222 => x"13050a00",
        2223 => x"97000000",
        2224 => x"e7000000",
        2225 => x"93090500",
        2226 => x"e31455fb",
        2227 => x"8357c900",
        2228 => x"93f70704",
        2229 => x"e39e07d0",
        2230 => x"03254102",
        2231 => x"6ff09fd1",
        2232 => x"b7260000",
        2233 => x"1307c100",
        2234 => x"9386c6e0",
        2235 => x"13060900",
        2236 => x"93050101",
        2237 => x"13050a00",
        2238 => x"ef00c01b",
        2239 => x"6ff09ffc",
        2240 => x"130101fd",
        2241 => x"232a5101",
        2242 => x"83a70501",
        2243 => x"930a0700",
        2244 => x"03a78500",
        2245 => x"23248102",
        2246 => x"23202103",
        2247 => x"232e3101",
        2248 => x"232c4101",
        2249 => x"23261102",
        2250 => x"23229102",
        2251 => x"23286101",
        2252 => x"23267101",
        2253 => x"93090500",
        2254 => x"13840500",
        2255 => x"13090600",
        2256 => x"138a0600",
        2257 => x"63d4e700",
        2258 => x"93070700",
        2259 => x"2320f900",
        2260 => x"03473404",
        2261 => x"63060700",
        2262 => x"93871700",
        2263 => x"2320f900",
        2264 => x"83270400",
        2265 => x"93f70702",
        2266 => x"63880700",
        2267 => x"83270900",
        2268 => x"93872700",
        2269 => x"2320f900",
        2270 => x"83240400",
        2271 => x"93f46400",
        2272 => x"639e0400",
        2273 => x"130b9401",
        2274 => x"930bf0ff",
        2275 => x"8327c400",
        2276 => x"03270900",
        2277 => x"b387e740",
        2278 => x"63c4f408",
        2279 => x"83473404",
        2280 => x"b336f000",
        2281 => x"83270400",
        2282 => x"93f70702",
        2283 => x"6392070c",
        2284 => x"13063404",
        2285 => x"93050a00",
        2286 => x"13850900",
        2287 => x"e7800a00",
        2288 => x"9307f0ff",
        2289 => x"630af506",
        2290 => x"83270400",
        2291 => x"13074000",
        2292 => x"93040000",
        2293 => x"93f76700",
        2294 => x"639ee700",
        2295 => x"83270900",
        2296 => x"8324c400",
        2297 => x"b384f440",
        2298 => x"93c7f4ff",
        2299 => x"93d7f741",
        2300 => x"b3f4f400",
        2301 => x"83278400",
        2302 => x"03270401",
        2303 => x"6356f700",
        2304 => x"b387e740",
        2305 => x"b384f400",
        2306 => x"13090000",
        2307 => x"1304a401",
        2308 => x"130bf0ff",
        2309 => x"63902409",
        2310 => x"13050000",
        2311 => x"6f000002",
        2312 => x"93061000",
        2313 => x"13060b00",
        2314 => x"93050a00",
        2315 => x"13850900",
        2316 => x"e7800a00",
        2317 => x"631a7503",
        2318 => x"1305f0ff",
        2319 => x"8320c102",
        2320 => x"03248102",
        2321 => x"83244102",
        2322 => x"03290102",
        2323 => x"8329c101",
        2324 => x"032a8101",
        2325 => x"832a4101",
        2326 => x"032b0101",
        2327 => x"832bc100",
        2328 => x"13010103",
        2329 => x"67800000",
        2330 => x"93841400",
        2331 => x"6ff01ff2",
        2332 => x"3307d400",
        2333 => x"13060003",
        2334 => x"a301c704",
        2335 => x"03475404",
        2336 => x"93871600",
        2337 => x"b307f400",
        2338 => x"93862600",
        2339 => x"a381e704",
        2340 => x"6ff01ff2",
        2341 => x"93061000",
        2342 => x"13060400",
        2343 => x"93050a00",
        2344 => x"13850900",
        2345 => x"e7800a00",
        2346 => x"e30865f9",
        2347 => x"13091900",
        2348 => x"6ff05ff6",
        2349 => x"130101fd",
        2350 => x"23248102",
        2351 => x"23229102",
        2352 => x"23202103",
        2353 => x"232e3101",
        2354 => x"23261102",
        2355 => x"232c4101",
        2356 => x"232a5101",
        2357 => x"23286101",
        2358 => x"83c88501",
        2359 => x"93078007",
        2360 => x"93040500",
        2361 => x"13840500",
        2362 => x"13090600",
        2363 => x"93890600",
        2364 => x"63ee1701",
        2365 => x"93072006",
        2366 => x"93863504",
        2367 => x"63ee1701",
        2368 => x"63840828",
        2369 => x"93078005",
        2370 => x"6380f822",
        2371 => x"930a2404",
        2372 => x"23011405",
        2373 => x"6f004004",
        2374 => x"9387d8f9",
        2375 => x"93f7f70f",
        2376 => x"13065001",
        2377 => x"e364f6fe",
        2378 => x"37360000",
        2379 => x"93972700",
        2380 => x"130606e0",
        2381 => x"b387c700",
        2382 => x"83a70700",
        2383 => x"67800700",
        2384 => x"83270700",
        2385 => x"938a2504",
        2386 => x"93864700",
        2387 => x"83a70700",
        2388 => x"2320d700",
        2389 => x"2381f504",
        2390 => x"93071000",
        2391 => x"6f008026",
        2392 => x"83a70500",
        2393 => x"03250700",
        2394 => x"13f60708",
        2395 => x"93054500",
        2396 => x"63060602",
        2397 => x"83270500",
        2398 => x"2320b700",
        2399 => x"37380000",
        2400 => x"63d80700",
        2401 => x"1307d002",
        2402 => x"b307f040",
        2403 => x"a301e404",
        2404 => x"130888dd",
        2405 => x"9308a000",
        2406 => x"6f004006",
        2407 => x"13f60704",
        2408 => x"83270500",
        2409 => x"2320b700",
        2410 => x"e30a06fc",
        2411 => x"93970701",
        2412 => x"93d70741",
        2413 => x"6ff09ffc",
        2414 => x"83a50500",
        2415 => x"03260700",
        2416 => x"13f50508",
        2417 => x"83270600",
        2418 => x"13064600",
        2419 => x"631a0500",
        2420 => x"93f50504",
        2421 => x"63860500",
        2422 => x"93970701",
        2423 => x"93d70701",
        2424 => x"2320c700",
        2425 => x"37380000",
        2426 => x"1307f006",
        2427 => x"130888dd",
        2428 => x"639ae814",
        2429 => x"93088000",
        2430 => x"a3010404",
        2431 => x"03274400",
        2432 => x"2324e400",
        2433 => x"634e0700",
        2434 => x"03260400",
        2435 => x"33e7e700",
        2436 => x"938a0600",
        2437 => x"1376b6ff",
        2438 => x"2320c400",
        2439 => x"63040702",
        2440 => x"938a0600",
        2441 => x"33f71703",
        2442 => x"938afaff",
        2443 => x"3307e800",
        2444 => x"03470700",
        2445 => x"2380ea00",
        2446 => x"13870700",
        2447 => x"b3d71703",
        2448 => x"e37217ff",
        2449 => x"93078000",
        2450 => x"6394f802",
        2451 => x"83270400",
        2452 => x"93f71700",
        2453 => x"638e0700",
        2454 => x"03274400",
        2455 => x"83270401",
        2456 => x"63c8e700",
        2457 => x"93070003",
        2458 => x"a38ffafe",
        2459 => x"938afaff",
        2460 => x"b3865641",
        2461 => x"2328d400",
        2462 => x"13870900",
        2463 => x"93060900",
        2464 => x"1306c100",
        2465 => x"93050400",
        2466 => x"13850400",
        2467 => x"eff05fc7",
        2468 => x"130af0ff",
        2469 => x"631e4513",
        2470 => x"1305f0ff",
        2471 => x"8320c102",
        2472 => x"03248102",
        2473 => x"83244102",
        2474 => x"03290102",
        2475 => x"8329c101",
        2476 => x"032a8101",
        2477 => x"832a4101",
        2478 => x"032b0101",
        2479 => x"13010103",
        2480 => x"67800000",
        2481 => x"83a70500",
        2482 => x"93e70702",
        2483 => x"23a0f500",
        2484 => x"37380000",
        2485 => x"93088007",
        2486 => x"1308c8de",
        2487 => x"a3021405",
        2488 => x"03260400",
        2489 => x"83250700",
        2490 => x"13750608",
        2491 => x"83a70500",
        2492 => x"93854500",
        2493 => x"631a0500",
        2494 => x"13750604",
        2495 => x"63060500",
        2496 => x"93970701",
        2497 => x"93d70701",
        2498 => x"2320b700",
        2499 => x"13771600",
        2500 => x"63060700",
        2501 => x"13660602",
        2502 => x"2320c400",
        2503 => x"638c0700",
        2504 => x"93080001",
        2505 => x"6ff05fed",
        2506 => x"37380000",
        2507 => x"130888dd",
        2508 => x"6ff0dffa",
        2509 => x"03270400",
        2510 => x"1377f7fd",
        2511 => x"2320e400",
        2512 => x"6ff01ffe",
        2513 => x"9308a000",
        2514 => x"6ff01feb",
        2515 => x"03a60500",
        2516 => x"83270700",
        2517 => x"83a54501",
        2518 => x"13780608",
        2519 => x"13854700",
        2520 => x"630a0800",
        2521 => x"2320a700",
        2522 => x"83a70700",
        2523 => x"23a0b700",
        2524 => x"6f008001",
        2525 => x"2320a700",
        2526 => x"13760604",
        2527 => x"83a70700",
        2528 => x"e30606fe",
        2529 => x"2390b700",
        2530 => x"23280400",
        2531 => x"938a0600",
        2532 => x"6ff09fee",
        2533 => x"83270700",
        2534 => x"03a64500",
        2535 => x"93050000",
        2536 => x"93864700",
        2537 => x"2320d700",
        2538 => x"83aa0700",
        2539 => x"13850a00",
        2540 => x"ef004009",
        2541 => x"63060500",
        2542 => x"33055541",
        2543 => x"2322a400",
        2544 => x"83274400",
        2545 => x"2328f400",
        2546 => x"a3010404",
        2547 => x"6ff0dfea",
        2548 => x"83260401",
        2549 => x"13860a00",
        2550 => x"93050900",
        2551 => x"13850400",
        2552 => x"e7800900",
        2553 => x"e30a45eb",
        2554 => x"83270400",
        2555 => x"93f72700",
        2556 => x"63940704",
        2557 => x"8327c100",
        2558 => x"0325c400",
        2559 => x"e350f5ea",
        2560 => x"13850700",
        2561 => x"6ff09fe9",
        2562 => x"93061000",
        2563 => x"13060b00",
        2564 => x"93050900",
        2565 => x"13850400",
        2566 => x"e7800900",
        2567 => x"e30e45e7",
        2568 => x"938a1a00",
        2569 => x"8327c400",
        2570 => x"0327c100",
        2571 => x"b387e740",
        2572 => x"e3ccfafc",
        2573 => x"6ff01ffc",
        2574 => x"930a0000",
        2575 => x"130b9401",
        2576 => x"6ff05ffe",
        2577 => x"93f5f50f",
        2578 => x"3306c500",
        2579 => x"6316c500",
        2580 => x"13050000",
        2581 => x"67800000",
        2582 => x"83470500",
        2583 => x"e38cb7fe",
        2584 => x"13051500",
        2585 => x"6ff09ffe",
        2586 => x"130101ff",
        2587 => x"23248100",
        2588 => x"23229100",
        2589 => x"13040500",
        2590 => x"13850500",
        2591 => x"93050600",
        2592 => x"23261100",
        2593 => x"23a80186",
        2594 => x"efe01fb7",
        2595 => x"9307f0ff",
        2596 => x"6318f500",
        2597 => x"83a70187",
        2598 => x"63840700",
        2599 => x"2320f400",
        2600 => x"8320c100",
        2601 => x"03248100",
        2602 => x"83244100",
        2603 => x"13010101",
        2604 => x"67800000",
        2605 => x"130101ff",
        2606 => x"23248100",
        2607 => x"23229100",
        2608 => x"13040500",
        2609 => x"13850500",
        2610 => x"23261100",
        2611 => x"23a80186",
        2612 => x"efe05fbb",
        2613 => x"9307f0ff",
        2614 => x"6318f500",
        2615 => x"83a70187",
        2616 => x"63840700",
        2617 => x"2320f400",
        2618 => x"8320c100",
        2619 => x"03248100",
        2620 => x"83244100",
        2621 => x"13010101",
        2622 => x"67800000",
        2623 => x"130101fe",
        2624 => x"232c8100",
        2625 => x"232e1100",
        2626 => x"232a9100",
        2627 => x"23282101",
        2628 => x"23263101",
        2629 => x"23244101",
        2630 => x"13040600",
        2631 => x"63940502",
        2632 => x"03248101",
        2633 => x"8320c101",
        2634 => x"83244101",
        2635 => x"03290101",
        2636 => x"8329c100",
        2637 => x"032a8100",
        2638 => x"93050600",
        2639 => x"13010102",
        2640 => x"6ff08fb0",
        2641 => x"63180602",
        2642 => x"eff04f98",
        2643 => x"93040000",
        2644 => x"8320c101",
        2645 => x"03248101",
        2646 => x"03290101",
        2647 => x"8329c100",
        2648 => x"032a8100",
        2649 => x"13850400",
        2650 => x"83244101",
        2651 => x"13010102",
        2652 => x"67800000",
        2653 => x"130a0500",
        2654 => x"93840500",
        2655 => x"ef008005",
        2656 => x"13090500",
        2657 => x"63668500",
        2658 => x"93571500",
        2659 => x"e3e287fc",
        2660 => x"93050400",
        2661 => x"13050a00",
        2662 => x"eff00fab",
        2663 => x"93090500",
        2664 => x"63160500",
        2665 => x"93840900",
        2666 => x"6ff09ffa",
        2667 => x"13060400",
        2668 => x"63748900",
        2669 => x"13060900",
        2670 => x"93850400",
        2671 => x"13850900",
        2672 => x"efe05f9d",
        2673 => x"93850400",
        2674 => x"13050a00",
        2675 => x"eff00f90",
        2676 => x"6ff05ffd",
        2677 => x"83a7c5ff",
        2678 => x"1385c7ff",
        2679 => x"63d80700",
        2680 => x"b385a500",
        2681 => x"83a70500",
        2682 => x"3305f500",
        2683 => x"67800000",
        2684 => x"30313233",
        2685 => x"34353637",
        2686 => x"38396162",
        2687 => x"63646566",
        2688 => x"00000000",
        2689 => x"a0040000",
        2690 => x"d8030000",
        2691 => x"d8030000",
        2692 => x"d8030000",
        2693 => x"ac040000",
        2694 => x"d8030000",
        2695 => x"d8030000",
        2696 => x"d8030000",
        2697 => x"d8030000",
        2698 => x"d8030000",
        2699 => x"d8030000",
        2700 => x"d8030000",
        2701 => x"d8030000",
        2702 => x"d8030000",
        2703 => x"d8030000",
        2704 => x"b8040000",
        2705 => x"d8030000",
        2706 => x"c4040000",
        2707 => x"d0040000",
        2708 => x"d8030000",
        2709 => x"dc040000",
        2710 => x"e8040000",
        2711 => x"d8030000",
        2712 => x"f4040000",
        2713 => x"94040000",
        2714 => x"d8030000",
        2715 => x"d8030000",
        2716 => x"d8030000",
        2717 => x"00050000",
        2718 => x"d8030000",
        2719 => x"d8030000",
        2720 => x"d8030000",
        2721 => x"d8030000",
        2722 => x"d8030000",
        2723 => x"d8030000",
        2724 => x"d8030000",
        2725 => x"10050000",
        2726 => x"a4050000",
        2727 => x"bc050000",
        2728 => x"ec050000",
        2729 => x"6c050000",
        2730 => x"6c050000",
        2731 => x"6c050000",
        2732 => x"6c050000",
        2733 => x"6c050000",
        2734 => x"6c050000",
        2735 => x"d4050000",
        2736 => x"6c050000",
        2737 => x"6c050000",
        2738 => x"6c050000",
        2739 => x"6c050000",
        2740 => x"84050000",
        2741 => x"84050000",
        2742 => x"a4050000",
        2743 => x"6c050000",
        2744 => x"6c050000",
        2745 => x"6c050000",
        2746 => x"6c050000",
        2747 => x"98050000",
        2748 => x"04060000",
        2749 => x"2c060000",
        2750 => x"6c050000",
        2751 => x"6c050000",
        2752 => x"6c050000",
        2753 => x"6c050000",
        2754 => x"6c050000",
        2755 => x"6c050000",
        2756 => x"6c050000",
        2757 => x"6c050000",
        2758 => x"6c050000",
        2759 => x"6c050000",
        2760 => x"6c050000",
        2761 => x"6c050000",
        2762 => x"6c050000",
        2763 => x"6c050000",
        2764 => x"84050000",
        2765 => x"84050000",
        2766 => x"6c050000",
        2767 => x"6c050000",
        2768 => x"6c050000",
        2769 => x"6c050000",
        2770 => x"6c050000",
        2771 => x"6c050000",
        2772 => x"6c050000",
        2773 => x"6c050000",
        2774 => x"6c050000",
        2775 => x"6c050000",
        2776 => x"6c050000",
        2777 => x"6c050000",
        2778 => x"98050000",
        2779 => x"00010202",
        2780 => x"03030303",
        2781 => x"04040404",
        2782 => x"04040404",
        2783 => x"05050505",
        2784 => x"05050505",
        2785 => x"05050505",
        2786 => x"05050505",
        2787 => x"06060606",
        2788 => x"06060606",
        2789 => x"06060606",
        2790 => x"06060606",
        2791 => x"06060606",
        2792 => x"06060606",
        2793 => x"06060606",
        2794 => x"06060606",
        2795 => x"07070707",
        2796 => x"07070707",
        2797 => x"07070707",
        2798 => x"07070707",
        2799 => x"07070707",
        2800 => x"07070707",
        2801 => x"07070707",
        2802 => x"07070707",
        2803 => x"07070707",
        2804 => x"07070707",
        2805 => x"07070707",
        2806 => x"07070707",
        2807 => x"07070707",
        2808 => x"07070707",
        2809 => x"07070707",
        2810 => x"07070707",
        2811 => x"08080808",
        2812 => x"08080808",
        2813 => x"08080808",
        2814 => x"08080808",
        2815 => x"08080808",
        2816 => x"08080808",
        2817 => x"08080808",
        2818 => x"08080808",
        2819 => x"08080808",
        2820 => x"08080808",
        2821 => x"08080808",
        2822 => x"08080808",
        2823 => x"08080808",
        2824 => x"08080808",
        2825 => x"08080808",
        2826 => x"08080808",
        2827 => x"08080808",
        2828 => x"08080808",
        2829 => x"08080808",
        2830 => x"08080808",
        2831 => x"08080808",
        2832 => x"08080808",
        2833 => x"08080808",
        2834 => x"08080808",
        2835 => x"08080808",
        2836 => x"08080808",
        2837 => x"08080808",
        2838 => x"08080808",
        2839 => x"08080808",
        2840 => x"08080808",
        2841 => x"08080808",
        2842 => x"08080808",
        2843 => x"0d0a4542",
        2844 => x"5245414b",
        2845 => x"21206d65",
        2846 => x"7063203d",
        2847 => x"20000000",
        2848 => x"20696e73",
        2849 => x"6e203d20",
        2850 => x"00000000",
        2851 => x"0d0a0000",
        2852 => x"0d0a0a44",
        2853 => x"6973706c",
        2854 => x"6179696e",
        2855 => x"67207468",
        2856 => x"65207469",
        2857 => x"6d652070",
        2858 => x"61737365",
        2859 => x"64207369",
        2860 => x"6e636520",
        2861 => x"72657365",
        2862 => x"740d0a0a",
        2863 => x"00000000",
        2864 => x"4f6e2d63",
        2865 => x"68697020",
        2866 => x"64656275",
        2867 => x"67676572",
        2868 => x"20666f75",
        2869 => x"6e642c20",
        2870 => x"736b6970",
        2871 => x"70696e67",
        2872 => x"20454252",
        2873 => x"45414b20",
        2874 => x"696e7374",
        2875 => x"72756374",
        2876 => x"696f6e0d",
        2877 => x"0a0d0a00",
        2878 => x"2530356c",
        2879 => x"643a2530",
        2880 => x"366c6420",
        2881 => x"20202530",
        2882 => x"326c643a",
        2883 => x"2530326c",
        2884 => x"643a2530",
        2885 => x"326c640d",
        2886 => x"00000000",
        2887 => x"696e7465",
        2888 => x"72727570",
        2889 => x"745f6469",
        2890 => x"72656374",
        2891 => x"00000000",
        2892 => x"54485541",
        2893 => x"53205249",
        2894 => x"53432d56",
        2895 => x"20525633",
        2896 => x"32494d20",
        2897 => x"62617265",
        2898 => x"206d6574",
        2899 => x"616c2070",
        2900 => x"726f6365",
        2901 => x"73736f72",
        2902 => x"00000000",
        2903 => x"54686520",
        2904 => x"48616775",
        2905 => x"6520556e",
        2906 => x"69766572",
        2907 => x"73697479",
        2908 => x"206f6620",
        2909 => x"4170706c",
        2910 => x"69656420",
        2911 => x"53636965",
        2912 => x"6e636573",
        2913 => x"00000000",
        2914 => x"44657061",
        2915 => x"72746d65",
        2916 => x"6e74206f",
        2917 => x"6620456c",
        2918 => x"65637472",
        2919 => x"6963616c",
        2920 => x"20456e67",
        2921 => x"696e6565",
        2922 => x"72696e67",
        2923 => x"00000000",
        2924 => x"4a2e452e",
        2925 => x"4a2e206f",
        2926 => x"70206465",
        2927 => x"6e204272",
        2928 => x"6f757700",
        2929 => x"232d302b",
        2930 => x"20000000",
        2931 => x"686c4c00",
        2932 => x"65666745",
        2933 => x"46470000",
        2934 => x"30313233",
        2935 => x"34353637",
        2936 => x"38394142",
        2937 => x"43444546",
        2938 => x"00000000",
        2939 => x"30313233",
        2940 => x"34353637",
        2941 => x"38396162",
        2942 => x"63646566",
        2943 => x"00000000",
        2944 => x"40250000",
        2945 => x"60250000",
        2946 => x"0c250000",
        2947 => x"0c250000",
        2948 => x"0c250000",
        2949 => x"0c250000",
        2950 => x"60250000",
        2951 => x"0c250000",
        2952 => x"0c250000",
        2953 => x"0c250000",
        2954 => x"0c250000",
        2955 => x"4c270000",
        2956 => x"b8250000",
        2957 => x"c4260000",
        2958 => x"0c250000",
        2959 => x"0c250000",
        2960 => x"94270000",
        2961 => x"0c250000",
        2962 => x"b8250000",
        2963 => x"0c250000",
        2964 => x"0c250000",
        2965 => x"d0260000",
        2966 => x"1c2d0000",
        2967 => x"302d0000",
        2968 => x"5c2d0000",
        2969 => x"882d0000",
        2970 => x"b02d0000",
        2971 => x"00000000",
        2972 => x"00000000",
        2973 => x"7c000020",
        2974 => x"e4000020",
        2975 => x"4c010020",
        2976 => x"00000000",
        2977 => x"00000000",
        2978 => x"00000000",
        2979 => x"00000000",
        2980 => x"00000000",
        2981 => x"00000000",
        2982 => x"00000000",
        2983 => x"00000000",
        2984 => x"00000000",
        2985 => x"00000000",
        2986 => x"00000000",
        2987 => x"00000000",
        2988 => x"00000000",
        2989 => x"00000000",
        2990 => x"00000000",
        2991 => x"18000020",
        2992 => x"00000000"
            );
end package rom_image;
