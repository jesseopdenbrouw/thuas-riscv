-- srec2vhdl table generator
-- for input file 'bootloader.srec'
-- date: Wed Nov 20 15:05:57 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package bootrom_image is
    constant bootrom_contents : memory_type := (
           0 => x"97020000",
           1 => x"93824262",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"37170010",
           8 => x"b7070020",
           9 => x"130747f6",
          10 => x"93870700",
          11 => x"37060020",
          12 => x"93060600",
          13 => x"63ecd70c",
          14 => x"b7070020",
          15 => x"93870700",
          16 => x"b7060020",
          17 => x"13870600",
          18 => x"63ece70c",
          19 => x"ef009030",
          20 => x"37c50100",
          21 => x"93051000",
          22 => x"13050520",
          23 => x"ef00c07c",
          24 => x"ef00902e",
          25 => x"37150010",
          26 => x"130545e0",
          27 => x"ef00d000",
          28 => x"732510fc",
          29 => x"37190010",
          30 => x"ef00d01b",
          31 => x"1305c9d7",
          32 => x"ef00807f",
          33 => x"370a00f0",
          34 => x"9307f03f",
          35 => x"93041000",
          36 => x"b709a000",
          37 => x"2322fa00",
          38 => x"b3899900",
          39 => x"9397c400",
          40 => x"639c0700",
          41 => x"1305a002",
          42 => x"ef00007b",
          43 => x"83274a00",
          44 => x"93d71700",
          45 => x"2322fa00",
          46 => x"ef000059",
          47 => x"13040500",
          48 => x"63160506",
          49 => x"93841400",
          50 => x"e39a34fd",
          51 => x"b70700f0",
          52 => x"23a20700",
          53 => x"631a0400",
          54 => x"93050000",
          55 => x"13050000",
          56 => x"ef008074",
          57 => x"e7000400",
          58 => x"ef000057",
          59 => x"1375f50f",
          60 => x"93071002",
          61 => x"6300f504",
          62 => x"93074002",
          63 => x"93040000",
          64 => x"6310f522",
          65 => x"13041000",
          66 => x"6f00c003",
          67 => x"83460700",
          68 => x"93871700",
          69 => x"13071700",
          70 => x"a38fd7fe",
          71 => x"6ff05ff1",
          72 => x"23800700",
          73 => x"93871700",
          74 => x"6ff0dff1",
          75 => x"13041000",
          76 => x"6ff0dff9",
          77 => x"37150010",
          78 => x"130585e3",
          79 => x"ef00c073",
          80 => x"13040000",
          81 => x"93040000",
          82 => x"b70900f0",
          83 => x"130b3005",
          84 => x"930ba004",
          85 => x"130c3002",
          86 => x"130a2000",
          87 => x"930ca000",
          88 => x"b71a0010",
          89 => x"83a74900",
          90 => x"93c71700",
          91 => x"23a2f900",
          92 => x"ef00804e",
          93 => x"1375f50f",
          94 => x"63186517",
          95 => x"ef00c04d",
          96 => x"137df50f",
          97 => x"9307fdfc",
          98 => x"93f7f70f",
          99 => x"6360fa10",
         100 => x"93071003",
         101 => x"6312fd04",
         102 => x"13052000",
         103 => x"ef00c071",
         104 => x"930dd5ff",
         105 => x"13054000",
         106 => x"ef000071",
         107 => x"130d0500",
         108 => x"b38dad00",
         109 => x"6318bd05",
         110 => x"130da000",
         111 => x"ef00c049",
         112 => x"1375f50f",
         113 => x"e31ca5ff",
         114 => x"e31e04f8",
         115 => x"13858ae3",
         116 => x"ef00806a",
         117 => x"6ff01ff9",
         118 => x"93072003",
         119 => x"13052000",
         120 => x"631afd00",
         121 => x"ef00406d",
         122 => x"930dc5ff",
         123 => x"13056000",
         124 => x"6ff09ffb",
         125 => x"ef00406c",
         126 => x"930db5ff",
         127 => x"13058000",
         128 => x"6ff09ffa",
         129 => x"1378cdff",
         130 => x"13052000",
         131 => x"23260101",
         132 => x"ef00806a",
         133 => x"0328c100",
         134 => x"93070500",
         135 => x"b70601ff",
         136 => x"37060001",
         137 => x"b705ffff",
         138 => x"13753d00",
         139 => x"93082000",
         140 => x"03270800",
         141 => x"9386f6ff",
         142 => x"13033000",
         143 => x"1306f6ff",
         144 => x"130e1000",
         145 => x"9385f50f",
         146 => x"63061503",
         147 => x"630a6502",
         148 => x"630cc501",
         149 => x"137707f0",
         150 => x"b3e7e700",
         151 => x"2320f800",
         152 => x"130d1d00",
         153 => x"6ff01ff5",
         154 => x"3377b700",
         155 => x"93978700",
         156 => x"6ff09ffe",
         157 => x"3377d700",
         158 => x"93970701",
         159 => x"6ff0dffd",
         160 => x"3377c700",
         161 => x"93978701",
         162 => x"6ff01ffd",
         163 => x"93079dfc",
         164 => x"93f7f70f",
         165 => x"6362fa04",
         166 => x"13052000",
         167 => x"ef00c061",
         168 => x"93077003",
         169 => x"13058000",
         170 => x"630afd00",
         171 => x"93078003",
         172 => x"13056000",
         173 => x"6304fd00",
         174 => x"13054000",
         175 => x"ef00c05f",
         176 => x"93040500",
         177 => x"130da000",
         178 => x"ef000039",
         179 => x"1375f50f",
         180 => x"e31ca5ff",
         181 => x"6ff05fef",
         182 => x"ef000038",
         183 => x"1375f50f",
         184 => x"e31c95ff",
         185 => x"6ff05fee",
         186 => x"631c7509",
         187 => x"63180400",
         188 => x"37150010",
         189 => x"130585e3",
         190 => x"ef000058",
         191 => x"93050000",
         192 => x"13050000",
         193 => x"ef004052",
         194 => x"b70700f0",
         195 => x"23a20700",
         196 => x"e7800400",
         197 => x"b70700f0",
         198 => x"1307a00a",
         199 => x"23a2e700",
         200 => x"97020000",
         201 => x"93824223",
         202 => x"73905230",
         203 => x"1305c9d7",
         204 => x"ef008054",
         205 => x"13040000",
         206 => x"b71a0010",
         207 => x"371b0010",
         208 => x"b7170010",
         209 => x"1385c7e3",
         210 => x"ef000053",
         211 => x"93059002",
         212 => x"13054101",
         213 => x"ef004032",
         214 => x"b7170010",
         215 => x"93090500",
         216 => x"938507e4",
         217 => x"13054101",
         218 => x"ef00002c",
         219 => x"631e0500",
         220 => x"37150010",
         221 => x"130545e4",
         222 => x"ef000050",
         223 => x"6f008003",
         224 => x"e31485e5",
         225 => x"6ff01ff9",
         226 => x"93850af3",
         227 => x"13054101",
         228 => x"ef008029",
         229 => x"63140502",
         230 => x"93050000",
         231 => x"ef00c048",
         232 => x"b70700f0",
         233 => x"23a20700",
         234 => x"93020000",
         235 => x"73905230",
         236 => x"e7800400",
         237 => x"e38609f8",
         238 => x"6f000019",
         239 => x"13063000",
         240 => x"93054bf3",
         241 => x"13054101",
         242 => x"ef009002",
         243 => x"63100504",
         244 => x"93050000",
         245 => x"13057101",
         246 => x"ef00405a",
         247 => x"93773500",
         248 => x"13040500",
         249 => x"63960706",
         250 => x"93058000",
         251 => x"ef00c06e",
         252 => x"37150010",
         253 => x"130585f3",
         254 => x"ef000048",
         255 => x"03250400",
         256 => x"93058000",
         257 => x"ef00406d",
         258 => x"6ff0dffa",
         259 => x"b7150010",
         260 => x"13063000",
         261 => x"938545f5",
         262 => x"13054101",
         263 => x"ef00407d",
         264 => x"631e0502",
         265 => x"93050101",
         266 => x"13057101",
         267 => x"ef000055",
         268 => x"93773500",
         269 => x"13040500",
         270 => x"639c0700",
         271 => x"03250101",
         272 => x"93050000",
         273 => x"ef008053",
         274 => x"2320a400",
         275 => x"6ff09ff6",
         276 => x"37150010",
         277 => x"1305c5f3",
         278 => x"6ff01ff2",
         279 => x"b7150010",
         280 => x"13063000",
         281 => x"938585f5",
         282 => x"13054101",
         283 => x"ef004078",
         284 => x"03474101",
         285 => x"9307e006",
         286 => x"6300050a",
         287 => x"631ef70a",
         288 => x"93773400",
         289 => x"e39607fc",
         290 => x"930b0404",
         291 => x"371c0010",
         292 => x"b71c0010",
         293 => x"371d0010",
         294 => x"930d80ff",
         295 => x"93058000",
         296 => x"13050400",
         297 => x"ef004063",
         298 => x"13058cf3",
         299 => x"ef00c03c",
         300 => x"83270400",
         301 => x"93058000",
         302 => x"93098001",
         303 => x"13850700",
         304 => x"2326f100",
         305 => x"ef004061",
         306 => x"1385ccf5",
         307 => x"ef00c03a",
         308 => x"370a00ff",
         309 => x"8327c100",
         310 => x"93069dc7",
         311 => x"33f54701",
         312 => x"33553501",
         313 => x"b306d500",
         314 => x"83c60600",
         315 => x"93f67609",
         316 => x"63800604",
         317 => x"938989ff",
         318 => x"ef000036",
         319 => x"135a8a00",
         320 => x"e39ab9fd",
         321 => x"13044400",
         322 => x"1305c9d7",
         323 => x"ef00c036",
         324 => x"e31674f9",
         325 => x"6ff0dfe2",
         326 => x"e304f7f6",
         327 => x"93050000",
         328 => x"13057101",
         329 => x"ef008045",
         330 => x"13040500",
         331 => x"6ff05ff5",
         332 => x"1305e002",
         333 => x"6ff01ffc",
         334 => x"e38409e0",
         335 => x"37150010",
         336 => x"130505f6",
         337 => x"ef004033",
         338 => x"1305c9d7",
         339 => x"ef00c032",
         340 => x"6ff01fdf",
         341 => x"130101fb",
         342 => x"23261104",
         343 => x"23245104",
         344 => x"23226104",
         345 => x"23207104",
         346 => x"232e8102",
         347 => x"232c9102",
         348 => x"232aa102",
         349 => x"2328b102",
         350 => x"2326c102",
         351 => x"2324d102",
         352 => x"2322e102",
         353 => x"2320f102",
         354 => x"232e0101",
         355 => x"232c1101",
         356 => x"232ac101",
         357 => x"2328d101",
         358 => x"2326e101",
         359 => x"2324f101",
         360 => x"73241034",
         361 => x"f3242034",
         362 => x"37150010",
         363 => x"130505df",
         364 => x"ef00802c",
         365 => x"93058000",
         366 => x"13850400",
         367 => x"ef00c051",
         368 => x"37150010",
         369 => x"1305c5d7",
         370 => x"ef00002b",
         371 => x"13044400",
         372 => x"73101434",
         373 => x"0324c103",
         374 => x"8320c104",
         375 => x"83228104",
         376 => x"03234104",
         377 => x"83230104",
         378 => x"83248103",
         379 => x"03254103",
         380 => x"83250103",
         381 => x"0326c102",
         382 => x"83268102",
         383 => x"03274102",
         384 => x"83270102",
         385 => x"0328c101",
         386 => x"83288101",
         387 => x"032e4101",
         388 => x"832e0101",
         389 => x"032fc100",
         390 => x"832f8100",
         391 => x"13010105",
         392 => x"73002030",
         393 => x"6f000000",
         394 => x"03460500",
         395 => x"83c60500",
         396 => x"13051500",
         397 => x"93851500",
         398 => x"6314d600",
         399 => x"e31606fe",
         400 => x"3305d640",
         401 => x"67800000",
         402 => x"b70700f0",
         403 => x"03a54710",
         404 => x"13758500",
         405 => x"67800000",
         406 => x"370700f0",
         407 => x"13070710",
         408 => x"83274700",
         409 => x"93f78700",
         410 => x"e38c07fe",
         411 => x"03258700",
         412 => x"1375f50f",
         413 => x"67800000",
         414 => x"130101fd",
         415 => x"232e3101",
         416 => x"b7190010",
         417 => x"23248102",
         418 => x"23229102",
         419 => x"23202103",
         420 => x"232c4101",
         421 => x"232a5101",
         422 => x"23286101",
         423 => x"23267101",
         424 => x"23261102",
         425 => x"93040500",
         426 => x"138bf5ff",
         427 => x"9389c9c2",
         428 => x"13040000",
         429 => x"13095001",
         430 => x"130a2000",
         431 => x"930a2001",
         432 => x"b71b0010",
         433 => x"eff05ff9",
         434 => x"1377f50f",
         435 => x"6340e902",
         436 => x"6352ea02",
         437 => x"9307d7ff",
         438 => x"63eefa00",
         439 => x"93972700",
         440 => x"b387f900",
         441 => x"83a70700",
         442 => x"67800700",
         443 => x"9307f007",
         444 => x"630cf706",
         445 => x"635c640f",
         446 => x"9377f50f",
         447 => x"938607fe",
         448 => x"93f6f60f",
         449 => x"1306e005",
         450 => x"e36ed6fa",
         451 => x"b3868400",
         452 => x"13050700",
         453 => x"2380f600",
         454 => x"13041400",
         455 => x"ef00c013",
         456 => x"6ff05ffa",
         457 => x"b3848400",
         458 => x"37150010",
         459 => x"23800400",
         460 => x"1305c5d7",
         461 => x"ef004014",
         462 => x"8320c102",
         463 => x"13050400",
         464 => x"03248102",
         465 => x"83244102",
         466 => x"03290102",
         467 => x"8329c101",
         468 => x"032a8101",
         469 => x"832a4101",
         470 => x"032b0101",
         471 => x"832bc100",
         472 => x"13010103",
         473 => x"67800000",
         474 => x"6354800a",
         475 => x"1305f007",
         476 => x"ef00800e",
         477 => x"1304f4ff",
         478 => x"6ff0dff4",
         479 => x"13850bd8",
         480 => x"ef00800f",
         481 => x"eff05fed",
         482 => x"1377f50f",
         483 => x"6346e902",
         484 => x"13040000",
         485 => x"6ff0dff3",
         486 => x"63508006",
         487 => x"1305f007",
         488 => x"1304f4ff",
         489 => x"ef00400b",
         490 => x"e31a04fe",
         491 => x"eff0dfea",
         492 => x"1377f50f",
         493 => x"e35ee9fc",
         494 => x"9307f007",
         495 => x"13040000",
         496 => x"e31af7f2",
         497 => x"23248101",
         498 => x"13040000",
         499 => x"130c5001",
         500 => x"13057000",
         501 => x"ef004008",
         502 => x"eff01fe8",
         503 => x"1377f50f",
         504 => x"634cec02",
         505 => x"032c8100",
         506 => x"6ff09fee",
         507 => x"13057000",
         508 => x"ef008006",
         509 => x"6ff01fed",
         510 => x"eff01fe6",
         511 => x"1377f50f",
         512 => x"93075001",
         513 => x"e3d6e7ec",
         514 => x"9307f007",
         515 => x"e314f7ee",
         516 => x"23248101",
         517 => x"6ff09ffb",
         518 => x"9307f007",
         519 => x"e30af7fa",
         520 => x"032c8100",
         521 => x"6ff01fed",
         522 => x"f32710fc",
         523 => x"63960700",
         524 => x"b7f7fa02",
         525 => x"93870708",
         526 => x"63060500",
         527 => x"33d5a702",
         528 => x"1305f5ff",
         529 => x"b70700f0",
         530 => x"23a6a710",
         531 => x"23a0b710",
         532 => x"23a20710",
         533 => x"67800000",
         534 => x"370700f0",
         535 => x"1375f50f",
         536 => x"13070710",
         537 => x"2324a700",
         538 => x"83274700",
         539 => x"93f70701",
         540 => x"e38c07fe",
         541 => x"67800000",
         542 => x"630e0502",
         543 => x"130101ff",
         544 => x"23248100",
         545 => x"23261100",
         546 => x"13040500",
         547 => x"03450500",
         548 => x"630a0500",
         549 => x"13041400",
         550 => x"eff01ffc",
         551 => x"03450400",
         552 => x"e31a05fe",
         553 => x"8320c100",
         554 => x"03248100",
         555 => x"13010101",
         556 => x"67800000",
         557 => x"67800000",
         558 => x"130101fe",
         559 => x"232e1100",
         560 => x"232c8100",
         561 => x"6350a00a",
         562 => x"23263101",
         563 => x"b7190010",
         564 => x"232a9100",
         565 => x"23282101",
         566 => x"23244101",
         567 => x"13090500",
         568 => x"938999c7",
         569 => x"93040000",
         570 => x"13040000",
         571 => x"130a1000",
         572 => x"6f000001",
         573 => x"3364c400",
         574 => x"93841400",
         575 => x"63029904",
         576 => x"eff09fd5",
         577 => x"b387a900",
         578 => x"83c70700",
         579 => x"130605fd",
         580 => x"13144400",
         581 => x"13f74700",
         582 => x"93f64704",
         583 => x"e31c07fc",
         584 => x"93f73700",
         585 => x"e38a06fc",
         586 => x"63944701",
         587 => x"13050502",
         588 => x"130595fa",
         589 => x"93841400",
         590 => x"3364a400",
         591 => x"e31299fc",
         592 => x"8320c101",
         593 => x"13050400",
         594 => x"03248101",
         595 => x"83244101",
         596 => x"03290101",
         597 => x"8329c100",
         598 => x"032a8100",
         599 => x"13010102",
         600 => x"67800000",
         601 => x"13040000",
         602 => x"8320c101",
         603 => x"13050400",
         604 => x"03248101",
         605 => x"13010102",
         606 => x"67800000",
         607 => x"83470500",
         608 => x"37160010",
         609 => x"130696c7",
         610 => x"3307f600",
         611 => x"03470700",
         612 => x"93060500",
         613 => x"13758700",
         614 => x"630e0500",
         615 => x"83c71600",
         616 => x"93861600",
         617 => x"3307f600",
         618 => x"03470700",
         619 => x"13758700",
         620 => x"e31605fe",
         621 => x"13754704",
         622 => x"630a0506",
         623 => x"13050000",
         624 => x"13031000",
         625 => x"6f000002",
         626 => x"83c71600",
         627 => x"93861600",
         628 => x"33e5a800",
         629 => x"3307f600",
         630 => x"03470700",
         631 => x"13784704",
         632 => x"63000804",
         633 => x"13784700",
         634 => x"938807fd",
         635 => x"13773700",
         636 => x"13154500",
         637 => x"e31a08fc",
         638 => x"63146700",
         639 => x"93870702",
         640 => x"938797fa",
         641 => x"93861600",
         642 => x"33e5a700",
         643 => x"83c70600",
         644 => x"3307f600",
         645 => x"03470700",
         646 => x"13784704",
         647 => x"e31408fc",
         648 => x"63840500",
         649 => x"23a0d500",
         650 => x"67800000",
         651 => x"13050000",
         652 => x"6ff01fff",
         653 => x"130101fe",
         654 => x"232e1100",
         655 => x"23220100",
         656 => x"23240100",
         657 => x"23260100",
         658 => x"630e0506",
         659 => x"232c8100",
         660 => x"13040500",
         661 => x"63400506",
         662 => x"b7d5cccc",
         663 => x"93064100",
         664 => x"9385d5cc",
         665 => x"13089000",
         666 => x"b337b402",
         667 => x"13060400",
         668 => x"13850600",
         669 => x"9386f6ff",
         670 => x"93d73700",
         671 => x"13972700",
         672 => x"3307f700",
         673 => x"13171700",
         674 => x"3304e440",
         675 => x"13040403",
         676 => x"a3858600",
         677 => x"13840700",
         678 => x"e368c8fc",
         679 => x"1305a500",
         680 => x"eff09fdd",
         681 => x"8320c101",
         682 => x"03248101",
         683 => x"13010102",
         684 => x"67800000",
         685 => x"1305d002",
         686 => x"eff01fda",
         687 => x"33048040",
         688 => x"6ff09ff9",
         689 => x"13050003",
         690 => x"eff01fd9",
         691 => x"8320c101",
         692 => x"13010102",
         693 => x"67800000",
         694 => x"130101fe",
         695 => x"232e1100",
         696 => x"23220100",
         697 => x"23240100",
         698 => x"23060100",
         699 => x"1387f5ff",
         700 => x"93077000",
         701 => x"93060500",
         702 => x"63e4e704",
         703 => x"93070700",
         704 => x"13054100",
         705 => x"b307f500",
         706 => x"b385b740",
         707 => x"13089003",
         708 => x"13f6f600",
         709 => x"13070603",
         710 => x"6374e800",
         711 => x"13077605",
         712 => x"2380e700",
         713 => x"9387f7ff",
         714 => x"93d64600",
         715 => x"e392f5fe",
         716 => x"eff09fd4",
         717 => x"8320c101",
         718 => x"13010102",
         719 => x"67800000",
         720 => x"93058000",
         721 => x"6ff0dffb",
         722 => x"37150010",
         723 => x"1305c5d8",
         724 => x"6ff09fd2",
         725 => x"130101ff",
         726 => x"23248100",
         727 => x"23229100",
         728 => x"37140010",
         729 => x"b7140010",
         730 => x"938744f6",
         731 => x"130444f6",
         732 => x"3304f440",
         733 => x"23202101",
         734 => x"23261100",
         735 => x"13542440",
         736 => x"938444f6",
         737 => x"13090000",
         738 => x"63108904",
         739 => x"b7140010",
         740 => x"37140010",
         741 => x"938744f6",
         742 => x"130444f6",
         743 => x"3304f440",
         744 => x"13542440",
         745 => x"938444f6",
         746 => x"13090000",
         747 => x"63188902",
         748 => x"8320c100",
         749 => x"03248100",
         750 => x"83244100",
         751 => x"03290100",
         752 => x"13010101",
         753 => x"67800000",
         754 => x"83a70400",
         755 => x"13091900",
         756 => x"93844400",
         757 => x"e7800700",
         758 => x"6ff01ffb",
         759 => x"83a70400",
         760 => x"13091900",
         761 => x"93844400",
         762 => x"e7800700",
         763 => x"6ff01ffc",
         764 => x"630a0602",
         765 => x"1306f6ff",
         766 => x"13070000",
         767 => x"b307e500",
         768 => x"b386e500",
         769 => x"83c70700",
         770 => x"83c60600",
         771 => x"6398d700",
         772 => x"6306c700",
         773 => x"13071700",
         774 => x"e39207fe",
         775 => x"3385d740",
         776 => x"67800000",
         777 => x"13050000",
         778 => x"67800000",
         779 => x"7c070010",
         780 => x"f4060010",
         781 => x"f4060010",
         782 => x"f4060010",
         783 => x"f4060010",
         784 => x"68070010",
         785 => x"f4060010",
         786 => x"24070010",
         787 => x"f4060010",
         788 => x"f4060010",
         789 => x"24070010",
         790 => x"f4060010",
         791 => x"f4060010",
         792 => x"f4060010",
         793 => x"f4060010",
         794 => x"f4060010",
         795 => x"f4060010",
         796 => x"f4060010",
         797 => x"98070010",
         798 => x"00202020",
         799 => x"20202020",
         800 => x"20202828",
         801 => x"28282820",
         802 => x"20202020",
         803 => x"20202020",
         804 => x"20202020",
         805 => x"20202020",
         806 => x"20881010",
         807 => x"10101010",
         808 => x"10101010",
         809 => x"10101010",
         810 => x"10040404",
         811 => x"04040404",
         812 => x"04040410",
         813 => x"10101010",
         814 => x"10104141",
         815 => x"41414141",
         816 => x"01010101",
         817 => x"01010101",
         818 => x"01010101",
         819 => x"01010101",
         820 => x"01010101",
         821 => x"10101010",
         822 => x"10104242",
         823 => x"42424242",
         824 => x"02020202",
         825 => x"02020202",
         826 => x"02020202",
         827 => x"02020202",
         828 => x"02020202",
         829 => x"10101010",
         830 => x"20000000",
         831 => x"00000000",
         832 => x"00000000",
         833 => x"00000000",
         834 => x"00000000",
         835 => x"00000000",
         836 => x"00000000",
         837 => x"00000000",
         838 => x"00000000",
         839 => x"00000000",
         840 => x"00000000",
         841 => x"00000000",
         842 => x"00000000",
         843 => x"00000000",
         844 => x"00000000",
         845 => x"00000000",
         846 => x"00000000",
         847 => x"00000000",
         848 => x"00000000",
         849 => x"00000000",
         850 => x"00000000",
         851 => x"00000000",
         852 => x"00000000",
         853 => x"00000000",
         854 => x"00000000",
         855 => x"00000000",
         856 => x"00000000",
         857 => x"00000000",
         858 => x"00000000",
         859 => x"00000000",
         860 => x"00000000",
         861 => x"00000000",
         862 => x"00000000",
         863 => x"0d0a0000",
         864 => x"3c627265",
         865 => x"616b3e0d",
         866 => x"0a000000",
         867 => x"0d0a5f5f",
         868 => x"5f202020",
         869 => x"20202020",
         870 => x"5f20205f",
         871 => x"5f202020",
         872 => x"205f205c",
         873 => x"202f5f5f",
         874 => x"205f5f20",
         875 => x"0d0a207c",
         876 => x"207c5f7c",
         877 => x"7c207c7c",
         878 => x"5f7c285f",
         879 => x"202d2d2d",
         880 => x"7c5f2920",
         881 => x"56205f5f",
         882 => x"29205f29",
         883 => x"0d0a207c",
         884 => x"207c207c",
         885 => x"7c5f7c7c",
         886 => x"207c5f5f",
         887 => x"29202020",
         888 => x"7c205c20",
         889 => x"20205f5f",
         890 => x"292f5f5f",
         891 => x"0d0a0000",
         892 => x"54726170",
         893 => x"3a206d63",
         894 => x"61757365",
         895 => x"203d2030",
         896 => x"78000000",
         897 => x"0d0a5448",
         898 => x"55415320",
         899 => x"52495343",
         900 => x"2d562042",
         901 => x"6f6f746c",
         902 => x"6f616465",
         903 => x"72207630",
         904 => x"2e362e33",
         905 => x"0d0a436c",
         906 => x"6f636b20",
         907 => x"66726571",
         908 => x"75656e63",
         909 => x"793a2000",
         910 => x"3f0a0000",
         911 => x"3e200000",
         912 => x"68000000",
         913 => x"48656c70",
         914 => x"3a0d0a20",
         915 => x"68202020",
         916 => x"20202020",
         917 => x"20202020",
         918 => x"20202020",
         919 => x"202d2074",
         920 => x"68697320",
         921 => x"68656c70",
         922 => x"0d0a2072",
         923 => x"20202020",
         924 => x"20202020",
         925 => x"20202020",
         926 => x"20202020",
         927 => x"2d207275",
         928 => x"6e206170",
         929 => x"706c6963",
         930 => x"6174696f",
         931 => x"6e0d0a20",
         932 => x"7277203c",
         933 => x"61646472",
         934 => x"3e202020",
         935 => x"20202020",
         936 => x"202d2072",
         937 => x"65616420",
         938 => x"776f7264",
         939 => x"2066726f",
         940 => x"6d206164",
         941 => x"64720d0a",
         942 => x"20777720",
         943 => x"3c616464",
         944 => x"723e203c",
         945 => x"64617461",
         946 => x"3e202d20",
         947 => x"77726974",
         948 => x"6520776f",
         949 => x"72642064",
         950 => x"61746120",
         951 => x"61742061",
         952 => x"6464720d",
         953 => x"0a206477",
         954 => x"203c6164",
         955 => x"64723e20",
         956 => x"20202020",
         957 => x"2020202d",
         958 => x"2064756d",
         959 => x"70203136",
         960 => x"20776f72",
         961 => x"64730d0a",
         962 => x"206e2020",
         963 => x"20202020",
         964 => x"20202020",
         965 => x"20202020",
         966 => x"20202d20",
         967 => x"64756d70",
         968 => x"206e6578",
         969 => x"74203136",
         970 => x"20776f72",
         971 => x"64730000",
         972 => x"72000000",
         973 => x"72772000",
         974 => x"3a200000",
         975 => x"4e6f7420",
         976 => x"6f6e2034",
         977 => x"2d627974",
         978 => x"6520626f",
         979 => x"756e6461",
         980 => x"72792100",
         981 => x"77772000",
         982 => x"64772000",
         983 => x"20200000",
         984 => x"3f3f0000",
         985 => x"00000000"
            );
end package bootrom_image;
