-- srec2vhdl table generator
-- for input file 'bootloader.srec'
-- date: Thu Jan  1 21:14:38 2026


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package bootrom_image is
    constant bootrom_contents : memory_type := (
           0 => x"97120000",
           1 => x"9382c28b",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"37060020",
           9 => x"13050500",
          10 => x"13060600",
          11 => x"637ac500",
          12 => x"b7150010",
          13 => x"3306a640",
          14 => x"9385c5fe",
          15 => x"ef00903f",
          16 => x"37050020",
          17 => x"37060020",
          18 => x"13050500",
          19 => x"13060600",
          20 => x"6378c500",
          21 => x"3306a640",
          22 => x"93050000",
          23 => x"ef00d03b",
          24 => x"37c50100",
          25 => x"93051000",
          26 => x"13050520",
          27 => x"ef005008",
          28 => x"ef00d039",
          29 => x"37150010",
          30 => x"130505cd",
          31 => x"ef00500c",
          32 => x"732530f1",
          33 => x"93058000",
          34 => x"ef005031",
          35 => x"37150010",
          36 => x"1305c5cf",
          37 => x"ef00d00a",
          38 => x"732510fc",
          39 => x"b71a0010",
          40 => x"ef005025",
          41 => x"13858acb",
          42 => x"ef009009",
          43 => x"b70900f0",
          44 => x"9307f03f",
          45 => x"3709a000",
          46 => x"23a2f900",
          47 => x"13091900",
          48 => x"93041000",
          49 => x"6f008001",
          50 => x"ef009001",
          51 => x"13040500",
          52 => x"93841400",
          53 => x"631a0502",
          54 => x"63822449",
          55 => x"9397c400",
          56 => x"e39407fe",
          57 => x"1305a002",
          58 => x"ef009003",
          59 => x"83a74900",
          60 => x"93841400",
          61 => x"93d71700",
          62 => x"23a2f900",
          63 => x"ef00407e",
          64 => x"13040500",
          65 => x"e30a05fc",
          66 => x"b70700f0",
          67 => x"23a20700",
          68 => x"ef00007b",
          69 => x"9377f50f",
          70 => x"13071002",
          71 => x"6380e762",
          72 => x"13074002",
          73 => x"6388e744",
          74 => x"23260100",
          75 => x"97020000",
          76 => x"9382c26b",
          77 => x"73905230",
          78 => x"371c0010",
          79 => x"13858acb",
          80 => x"ef001000",
          81 => x"130c4cd1",
          82 => x"13090000",
          83 => x"13045001",
          84 => x"930c7002",
          85 => x"9304a000",
          86 => x"13050c00",
          87 => x"ef00407e",
          88 => x"130b0000",
          89 => x"130af007",
          90 => x"9309d000",
          91 => x"ef004075",
          92 => x"13070500",
          93 => x"1375f50f",
          94 => x"630c8504",
          95 => x"6346a402",
          96 => x"63049506",
          97 => x"63023507",
          98 => x"93068000",
          99 => x"6300d502",
         100 => x"63d86c11",
         101 => x"ef00c072",
         102 => x"13070500",
         103 => x"1375f50f",
         104 => x"630a8502",
         105 => x"e35ea4fc",
         106 => x"e31445ff",
         107 => x"631c0b10",
         108 => x"ef000071",
         109 => x"13070500",
         110 => x"1375f50f",
         111 => x"e31085fc",
         112 => x"ef000070",
         113 => x"13070500",
         114 => x"1375f50f",
         115 => x"e31885fa",
         116 => x"630a0b28",
         117 => x"1305f007",
         118 => x"130bfbff",
         119 => x"ef004074",
         120 => x"e31a0bfe",
         121 => x"6ff09ff8",
         122 => x"b3072b00",
         123 => x"23820702",
         124 => x"13858acb",
         125 => x"ef00c074",
         126 => x"83574102",
         127 => x"13078006",
         128 => x"638ae70c",
         129 => x"13072007",
         130 => x"6380e70e",
         131 => x"37670000",
         132 => x"13072727",
         133 => x"6380e710",
         134 => x"03574102",
         135 => x"b7670000",
         136 => x"93877727",
         137 => x"630cf712",
         138 => x"03574102",
         139 => x"b7770000",
         140 => x"93872787",
         141 => x"630ef714",
         142 => x"03574102",
         143 => x"b7770000",
         144 => x"93877787",
         145 => x"630af718",
         146 => x"03574102",
         147 => x"b7770000",
         148 => x"93872777",
         149 => x"630cf71a",
         150 => x"03574102",
         151 => x"b7770000",
         152 => x"93877777",
         153 => x"630af720",
         154 => x"03574102",
         155 => x"b7770000",
         156 => x"93874776",
         157 => x"630cf722",
         158 => x"03574102",
         159 => x"9307e006",
         160 => x"630cf722",
         161 => x"e30a0bec",
         162 => x"b7170010",
         163 => x"138547ee",
         164 => x"ef00006b",
         165 => x"13858acb",
         166 => x"ef00806a",
         167 => x"6ff0dfeb",
         168 => x"930607fe",
         169 => x"93f6f60f",
         170 => x"1306e005",
         171 => x"e360d6ec",
         172 => x"b3062b00",
         173 => x"2382e602",
         174 => x"130b1b00",
         175 => x"ef004066",
         176 => x"6ff0dfea",
         177 => x"1305f007",
         178 => x"ef008065",
         179 => x"130bfbff",
         180 => x"6ff0dfe9",
         181 => x"b7170010",
         182 => x"1385c7d1",
         183 => x"ef004066",
         184 => x"e30c0be6",
         185 => x"6ff01ffb",
         186 => x"93050000",
         187 => x"13050000",
         188 => x"ef000060",
         189 => x"b70700f0",
         190 => x"23a20700",
         191 => x"93020000",
         192 => x"73905230",
         193 => x"8327c100",
         194 => x"e7800700",
         195 => x"e3060be4",
         196 => x"6ff05ff8",
         197 => x"03476102",
         198 => x"93070002",
         199 => x"e31ef7ee",
         200 => x"93050000",
         201 => x"13057102",
         202 => x"ef00c071",
         203 => x"93058000",
         204 => x"83490500",
         205 => x"13090500",
         206 => x"ef005006",
         207 => x"b7170010",
         208 => x"138587cf",
         209 => x"ef00c05f",
         210 => x"13850900",
         211 => x"93052000",
         212 => x"ef00d004",
         213 => x"e3020be0",
         214 => x"6ff0dff3",
         215 => x"03476102",
         216 => x"93070002",
         217 => x"e312f7ec",
         218 => x"b305e100",
         219 => x"13057102",
         220 => x"ef00406d",
         221 => x"13090500",
         222 => x"03250102",
         223 => x"93050000",
         224 => x"ef00406c",
         225 => x"2300a900",
         226 => x"e3080bdc",
         227 => x"6ff09ff0",
         228 => x"03476102",
         229 => x"93070002",
         230 => x"e310f7ea",
         231 => x"93050000",
         232 => x"13057102",
         233 => x"ef00006a",
         234 => x"93058000",
         235 => x"83590500",
         236 => x"13090500",
         237 => x"ef00807e",
         238 => x"b7170010",
         239 => x"138587cf",
         240 => x"ef000058",
         241 => x"13850900",
         242 => x"93054000",
         243 => x"ef00007d",
         244 => x"e3040bd8",
         245 => x"6ff01fec",
         246 => x"03476102",
         247 => x"93070002",
         248 => x"e314f7e6",
         249 => x"b305e100",
         250 => x"13057102",
         251 => x"ef008065",
         252 => x"13090500",
         253 => x"03250102",
         254 => x"93050000",
         255 => x"ef008064",
         256 => x"2310a900",
         257 => x"e30a0bd4",
         258 => x"6ff0dfe8",
         259 => x"03476102",
         260 => x"93070002",
         261 => x"e312f7e4",
         262 => x"93050000",
         263 => x"13057102",
         264 => x"ef004062",
         265 => x"93058000",
         266 => x"83290500",
         267 => x"13090500",
         268 => x"ef00c076",
         269 => x"b7170010",
         270 => x"138587cf",
         271 => x"ef004050",
         272 => x"13850900",
         273 => x"93058000",
         274 => x"ef004075",
         275 => x"e3060bd0",
         276 => x"6ff05fe4",
         277 => x"ef00c046",
         278 => x"13070500",
         279 => x"1375f50f",
         280 => x"e31e85d0",
         281 => x"ef00c045",
         282 => x"13070500",
         283 => x"1375f50f",
         284 => x"e31685d0",
         285 => x"6ff01ffe",
         286 => x"03476102",
         287 => x"93070002",
         288 => x"e314f7de",
         289 => x"b305e100",
         290 => x"13057102",
         291 => x"ef00805b",
         292 => x"13090500",
         293 => x"03250102",
         294 => x"93050000",
         295 => x"ef00805a",
         296 => x"2320a900",
         297 => x"e30a0bca",
         298 => x"6ff0dfde",
         299 => x"03476102",
         300 => x"93070002",
         301 => x"e312f7dc",
         302 => x"03474102",
         303 => x"9307e006",
         304 => x"630af700",
         305 => x"93050000",
         306 => x"13057102",
         307 => x"ef008057",
         308 => x"13090500",
         309 => x"137ac9ff",
         310 => x"13090a04",
         311 => x"930be005",
         312 => x"130b80ff",
         313 => x"93058000",
         314 => x"13050a00",
         315 => x"ef00006b",
         316 => x"b7170010",
         317 => x"138587cf",
         318 => x"ef008044",
         319 => x"83290a00",
         320 => x"93058000",
         321 => x"130d8001",
         322 => x"13850900",
         323 => x"ef000069",
         324 => x"b7170010",
         325 => x"138507ee",
         326 => x"ef008042",
         327 => x"b70d00ff",
         328 => x"33f5b901",
         329 => x"3355a501",
         330 => x"930605fe",
         331 => x"63f4db00",
         332 => x"1305e002",
         333 => x"130d8dff",
         334 => x"ef00803e",
         335 => x"93dd8d00",
         336 => x"e3106dff",
         337 => x"b7170010",
         338 => x"130a4a00",
         339 => x"138587cb",
         340 => x"ef00003f",
         341 => x"e3182af9",
         342 => x"6ff01fc0",
         343 => x"b70700f0",
         344 => x"23a20700",
         345 => x"93050000",
         346 => x"ef008038",
         347 => x"e7000400",
         348 => x"6ff01fba",
         349 => x"13091000",
         350 => x"371b0010",
         351 => x"93070bd1",
         352 => x"23260100",
         353 => x"b70400f0",
         354 => x"93093005",
         355 => x"130ca004",
         356 => x"930b3002",
         357 => x"930d2000",
         358 => x"130aa000",
         359 => x"232ef100",
         360 => x"83a74400",
         361 => x"93c71700",
         362 => x"23a2f400",
         363 => x"ef004031",
         364 => x"9377f50f",
         365 => x"63883703",
         366 => x"638e8705",
         367 => x"638c7707",
         368 => x"e31009fe",
         369 => x"0325c101",
         370 => x"ef008037",
         371 => x"83a74400",
         372 => x"93c71700",
         373 => x"23a2f400",
         374 => x"ef00802e",
         375 => x"9377f50f",
         376 => x"e39c37fd",
         377 => x"ef00c02d",
         378 => x"1374f50f",
         379 => x"9307f4fc",
         380 => x"93f7f70f",
         381 => x"63f6fd08",
         382 => x"930794fc",
         383 => x"93f7f70f",
         384 => x"63f2fd04",
         385 => x"ef00c02b",
         386 => x"9377f50f",
         387 => x"e39c47ff",
         388 => x"6ff01ffb",
         389 => x"63060914",
         390 => x"93050000",
         391 => x"13050000",
         392 => x"ef00002d",
         393 => x"b70700f0",
         394 => x"23a20700",
         395 => x"8327c100",
         396 => x"e7800700",
         397 => x"b70700f0",
         398 => x"1307a00a",
         399 => x"23a2e700",
         400 => x"6ff0dfae",
         401 => x"13052000",
         402 => x"ef008033",
         403 => x"93077003",
         404 => x"6304f418",
         405 => x"93078003",
         406 => x"630cf40e",
         407 => x"13054000",
         408 => x"ef000032",
         409 => x"13040500",
         410 => x"930ca000",
         411 => x"ef004025",
         412 => x"9377f50f",
         413 => x"e39c97ff",
         414 => x"23268100",
         415 => x"6ff05ff4",
         416 => x"93071003",
         417 => x"630af412",
         418 => x"93072003",
         419 => x"13052000",
         420 => x"630ef40c",
         421 => x"ef00c02e",
         422 => x"13040500",
         423 => x"13058000",
         424 => x"ef00002e",
         425 => x"1304b4ff",
         426 => x"930c0500",
         427 => x"630c040e",
         428 => x"b70701ff",
         429 => x"9387f7ff",
         430 => x"b7060001",
         431 => x"2328f100",
         432 => x"9387f6ff",
         433 => x"232af100",
         434 => x"b707ffff",
         435 => x"9387f70f",
         436 => x"33049401",
         437 => x"232cf100",
         438 => x"6f004003",
         439 => x"93073000",
         440 => x"6308f70a",
         441 => x"83278101",
         442 => x"13f806f0",
         443 => x"93158500",
         444 => x"b3f6f600",
         445 => x"93071000",
         446 => x"6308f708",
         447 => x"33670501",
         448 => x"2320ed00",
         449 => x"938c1c00",
         450 => x"638e8c08",
         451 => x"13052000",
         452 => x"ef000027",
         453 => x"13fdccff",
         454 => x"13f73c00",
         455 => x"93072000",
         456 => x"83260d00",
         457 => x"e31cf7fa",
         458 => x"83270101",
         459 => x"13170501",
         460 => x"b3f6f600",
         461 => x"3367d700",
         462 => x"6ff09ffc",
         463 => x"371b0010",
         464 => x"13050bd1",
         465 => x"ef00c01f",
         466 => x"13090000",
         467 => x"6ff01fe3",
         468 => x"13056000",
         469 => x"ef00c022",
         470 => x"13040500",
         471 => x"6ff0dff0",
         472 => x"13050bd1",
         473 => x"ef00c01d",
         474 => x"6ff01feb",
         475 => x"ef004021",
         476 => x"13040500",
         477 => x"13056000",
         478 => x"ef008020",
         479 => x"1304c4ff",
         480 => x"930c0500",
         481 => x"6ff09ff2",
         482 => x"33e7d500",
         483 => x"6ff05ff7",
         484 => x"83274101",
         485 => x"13178501",
         486 => x"b3f6f600",
         487 => x"3367d700",
         488 => x"6ff01ff6",
         489 => x"1304a000",
         490 => x"ef008011",
         491 => x"9377f50f",
         492 => x"e39c87fe",
         493 => x"6ff0dfe0",
         494 => x"13052000",
         495 => x"ef00401c",
         496 => x"13040500",
         497 => x"13054000",
         498 => x"ef00801b",
         499 => x"1304d4ff",
         500 => x"930c0500",
         501 => x"6ff09fed",
         502 => x"13058000",
         503 => x"ef00401a",
         504 => x"13040500",
         505 => x"6ff05fe8",
         506 => x"130101fb",
         507 => x"23261104",
         508 => x"23245104",
         509 => x"23226104",
         510 => x"23207104",
         511 => x"232e8102",
         512 => x"232c9102",
         513 => x"232aa102",
         514 => x"2328b102",
         515 => x"2326c102",
         516 => x"2324d102",
         517 => x"2322e102",
         518 => x"2320f102",
         519 => x"232e0101",
         520 => x"232c1101",
         521 => x"232ac101",
         522 => x"2328d101",
         523 => x"2326e101",
         524 => x"2324f101",
         525 => x"73241034",
         526 => x"f3242034",
         527 => x"37150010",
         528 => x"1305c5cb",
         529 => x"ef00c00f",
         530 => x"13850400",
         531 => x"93058000",
         532 => x"ef00c034",
         533 => x"37150010",
         534 => x"130585cb",
         535 => x"ef00400e",
         536 => x"63c40400",
         537 => x"13044400",
         538 => x"73101434",
         539 => x"0324c103",
         540 => x"8320c104",
         541 => x"83228104",
         542 => x"03234104",
         543 => x"83230104",
         544 => x"83248103",
         545 => x"03254103",
         546 => x"83250103",
         547 => x"0326c102",
         548 => x"83268102",
         549 => x"03274102",
         550 => x"83270102",
         551 => x"0328c101",
         552 => x"83288101",
         553 => x"032e4101",
         554 => x"832e0101",
         555 => x"032fc100",
         556 => x"832f8100",
         557 => x"13010105",
         558 => x"73002030",
         559 => x"6f000000",
         560 => x"370700f0",
         561 => x"13070710",
         562 => x"83274700",
         563 => x"93f78700",
         564 => x"e38c07fe",
         565 => x"03258700",
         566 => x"1375f50f",
         567 => x"67800000",
         568 => x"b70700f0",
         569 => x"03a54710",
         570 => x"13758500",
         571 => x"67800000",
         572 => x"f32710fc",
         573 => x"63960700",
         574 => x"b7f7fa02",
         575 => x"93870708",
         576 => x"63060500",
         577 => x"33d5a702",
         578 => x"1305f5ff",
         579 => x"b70700f0",
         580 => x"23a6a710",
         581 => x"23a0b710",
         582 => x"23a20710",
         583 => x"67800000",
         584 => x"370700f0",
         585 => x"1375f50f",
         586 => x"13070710",
         587 => x"2324a700",
         588 => x"83274700",
         589 => x"93f70701",
         590 => x"e38c07fe",
         591 => x"67800000",
         592 => x"630e0502",
         593 => x"130101ff",
         594 => x"23248100",
         595 => x"23261100",
         596 => x"13040500",
         597 => x"03450500",
         598 => x"630a0500",
         599 => x"13041400",
         600 => x"eff01ffc",
         601 => x"03450400",
         602 => x"e31a05fe",
         603 => x"8320c100",
         604 => x"03248100",
         605 => x"13010101",
         606 => x"67800000",
         607 => x"67800000",
         608 => x"130101fe",
         609 => x"232e1100",
         610 => x"232c8100",
         611 => x"6350a00a",
         612 => x"23263101",
         613 => x"b7190010",
         614 => x"232a9100",
         615 => x"23282101",
         616 => x"23244101",
         617 => x"13090500",
         618 => x"938999ee",
         619 => x"93040000",
         620 => x"13040000",
         621 => x"130a1000",
         622 => x"6f000001",
         623 => x"3364c400",
         624 => x"93841400",
         625 => x"63029904",
         626 => x"eff09fef",
         627 => x"b387a900",
         628 => x"83c70700",
         629 => x"130605fd",
         630 => x"13144400",
         631 => x"13f74700",
         632 => x"93f64704",
         633 => x"e31c07fc",
         634 => x"93f73700",
         635 => x"e38a06fc",
         636 => x"63944701",
         637 => x"13050502",
         638 => x"130595fa",
         639 => x"93841400",
         640 => x"3364a400",
         641 => x"e31299fc",
         642 => x"8320c101",
         643 => x"13050400",
         644 => x"03248101",
         645 => x"83244101",
         646 => x"03290101",
         647 => x"8329c100",
         648 => x"032a8100",
         649 => x"13010102",
         650 => x"67800000",
         651 => x"13040000",
         652 => x"8320c101",
         653 => x"13050400",
         654 => x"03248101",
         655 => x"13010102",
         656 => x"67800000",
         657 => x"83470500",
         658 => x"37160010",
         659 => x"130696ee",
         660 => x"3307f600",
         661 => x"03470700",
         662 => x"93060500",
         663 => x"13758700",
         664 => x"630e0500",
         665 => x"83c71600",
         666 => x"93861600",
         667 => x"3307f600",
         668 => x"03470700",
         669 => x"13758700",
         670 => x"e31605fe",
         671 => x"13754704",
         672 => x"63040506",
         673 => x"13050000",
         674 => x"13031000",
         675 => x"6f000002",
         676 => x"83c71600",
         677 => x"93861600",
         678 => x"33e5a800",
         679 => x"3307f600",
         680 => x"03470700",
         681 => x"13784704",
         682 => x"63000804",
         683 => x"13784700",
         684 => x"938807fd",
         685 => x"13773700",
         686 => x"13154500",
         687 => x"e31a08fc",
         688 => x"63146700",
         689 => x"93870702",
         690 => x"938797fa",
         691 => x"93861600",
         692 => x"33e5a700",
         693 => x"83c70600",
         694 => x"3307f600",
         695 => x"03470700",
         696 => x"13784704",
         697 => x"e31408fc",
         698 => x"63840500",
         699 => x"23a0d500",
         700 => x"67800000",
         701 => x"130101fd",
         702 => x"23261102",
         703 => x"232a0100",
         704 => x"232c0100",
         705 => x"232e0100",
         706 => x"63000508",
         707 => x"93070500",
         708 => x"63400506",
         709 => x"b7d5cccc",
         710 => x"13850700",
         711 => x"9385d5cc",
         712 => x"93064101",
         713 => x"93089000",
         714 => x"b337b502",
         715 => x"13060500",
         716 => x"13880600",
         717 => x"9386f6ff",
         718 => x"93d73700",
         719 => x"13972700",
         720 => x"3307f700",
         721 => x"13171700",
         722 => x"3305e540",
         723 => x"13050503",
         724 => x"a385a600",
         725 => x"13850700",
         726 => x"e3e8c8fc",
         727 => x"1305a800",
         728 => x"eff01fde",
         729 => x"8320c102",
         730 => x"13010103",
         731 => x"67800000",
         732 => x"2326a100",
         733 => x"1305d002",
         734 => x"eff09fda",
         735 => x"8327c100",
         736 => x"b307f040",
         737 => x"6ff01ff9",
         738 => x"13050003",
         739 => x"eff05fd9",
         740 => x"8320c102",
         741 => x"13010103",
         742 => x"67800000",
         743 => x"130101fe",
         744 => x"232e1100",
         745 => x"23220100",
         746 => x"23240100",
         747 => x"23060100",
         748 => x"1387f5ff",
         749 => x"93077000",
         750 => x"93060500",
         751 => x"63e4e704",
         752 => x"93070700",
         753 => x"13054100",
         754 => x"b307f500",
         755 => x"b385b740",
         756 => x"13089003",
         757 => x"13f6f600",
         758 => x"13070603",
         759 => x"6374e800",
         760 => x"13077605",
         761 => x"2380e700",
         762 => x"9387f7ff",
         763 => x"93d64600",
         764 => x"e392f5fe",
         765 => x"eff0dfd4",
         766 => x"8320c101",
         767 => x"13010102",
         768 => x"67800000",
         769 => x"93058000",
         770 => x"6ff0dffb",
         771 => x"37150010",
         772 => x"130585c5",
         773 => x"6ff0dfd2",
         774 => x"13030500",
         775 => x"630a0600",
         776 => x"2300b300",
         777 => x"1306f6ff",
         778 => x"13031300",
         779 => x"e31a06fe",
         780 => x"67800000",
         781 => x"13030500",
         782 => x"630e0600",
         783 => x"83830500",
         784 => x"23007300",
         785 => x"1306f6ff",
         786 => x"13031300",
         787 => x"93851500",
         788 => x"e31606fe",
         789 => x"67800000",
         790 => x"0d0a5f5f",
         791 => x"5f202020",
         792 => x"20202020",
         793 => x"5f20205f",
         794 => x"5f202020",
         795 => x"205f205c",
         796 => x"202f5f5f",
         797 => x"205f5f20",
         798 => x"0d0a207c",
         799 => x"207c5f7c",
         800 => x"7c207c7c",
         801 => x"5f7c285f",
         802 => x"202d2d2d",
         803 => x"7c5f2920",
         804 => x"56205f5f",
         805 => x"29205f29",
         806 => x"0d0a207c",
         807 => x"207c207c",
         808 => x"7c5f7c7c",
         809 => x"207c5f5f",
         810 => x"29202020",
         811 => x"7c205c20",
         812 => x"20205f5f",
         813 => x"292f5f5f",
         814 => x"0d0a0000",
         815 => x"54726170",
         816 => x"3a206d63",
         817 => x"61757365",
         818 => x"203d2030",
         819 => x"78000000",
         820 => x"0d0a5448",
         821 => x"55415320",
         822 => x"52495343",
         823 => x"2d562042",
         824 => x"6f6f746c",
         825 => x"6f616465",
         826 => x"72207630",
         827 => x"2e370d0a",
         828 => x"48617264",
         829 => x"77617265",
         830 => x"3a200000",
         831 => x"0d0a436c",
         832 => x"6f636b20",
         833 => x"66726571",
         834 => x"75656e63",
         835 => x"793a2000",
         836 => x"3f0a0000",
         837 => x"3e200000",
         838 => x"68000000",
         839 => x"48656c70",
         840 => x"3a0d0a20",
         841 => x"68202020",
         842 => x"20202020",
         843 => x"20202020",
         844 => x"20202020",
         845 => x"202d2074",
         846 => x"68697320",
         847 => x"68656c70",
         848 => x"0d0a2072",
         849 => x"20202020",
         850 => x"20202020",
         851 => x"20202020",
         852 => x"20202020",
         853 => x"2d207275",
         854 => x"6e206170",
         855 => x"706c6963",
         856 => x"6174696f",
         857 => x"6e0d0a20",
         858 => x"7262203c",
         859 => x"61646472",
         860 => x"3e202020",
         861 => x"20202020",
         862 => x"202d2072",
         863 => x"65616420",
         864 => x"62797465",
         865 => x"2066726f",
         866 => x"6d206164",
         867 => x"64720d0a",
         868 => x"20776220",
         869 => x"3c616464",
         870 => x"723e203c",
         871 => x"64617461",
         872 => x"3e202d20",
         873 => x"77726974",
         874 => x"65206279",
         875 => x"74652064",
         876 => x"61746120",
         877 => x"61742061",
         878 => x"6464720d",
         879 => x"0a207268",
         880 => x"203c6164",
         881 => x"64723e20",
         882 => x"20202020",
         883 => x"2020202d",
         884 => x"20726561",
         885 => x"64206861",
         886 => x"6c66776f",
         887 => x"72642066",
         888 => x"726f6d20",
         889 => x"61646472",
         890 => x"0d0a2077",
         891 => x"68203c61",
         892 => x"6464723e",
         893 => x"203c6461",
         894 => x"74613e20",
         895 => x"2d207772",
         896 => x"69746520",
         897 => x"68616c66",
         898 => x"776f7264",
         899 => x"20646174",
         900 => x"61206174",
         901 => x"20616464",
         902 => x"720d0a20",
         903 => x"7277203c",
         904 => x"61646472",
         905 => x"3e202020",
         906 => x"20202020",
         907 => x"202d2072",
         908 => x"65616420",
         909 => x"776f7264",
         910 => x"2066726f",
         911 => x"6d206164",
         912 => x"64720d0a",
         913 => x"20777720",
         914 => x"3c616464",
         915 => x"723e203c",
         916 => x"64617461",
         917 => x"3e202d20",
         918 => x"77726974",
         919 => x"6520776f",
         920 => x"72642064",
         921 => x"61746120",
         922 => x"61742061",
         923 => x"6464720d",
         924 => x"0a206477",
         925 => x"203c6164",
         926 => x"64723e20",
         927 => x"20202020",
         928 => x"2020202d",
         929 => x"2064756d",
         930 => x"70203136",
         931 => x"20776f72",
         932 => x"64730d0a",
         933 => x"206e2020",
         934 => x"20202020",
         935 => x"20202020",
         936 => x"20202020",
         937 => x"20202d20",
         938 => x"64756d70",
         939 => x"206e6578",
         940 => x"74203136",
         941 => x"20776f72",
         942 => x"64730000",
         943 => x"72000000",
         944 => x"72622000",
         945 => x"77622000",
         946 => x"72682000",
         947 => x"77682000",
         948 => x"72772000",
         949 => x"77772000",
         950 => x"64772000",
         951 => x"6e000000",
         952 => x"20200000",
         953 => x"3f3f0000",
         954 => x"00202020",
         955 => x"20202020",
         956 => x"20202828",
         957 => x"28282820",
         958 => x"20202020",
         959 => x"20202020",
         960 => x"20202020",
         961 => x"20202020",
         962 => x"20881010",
         963 => x"10101010",
         964 => x"10101010",
         965 => x"10101010",
         966 => x"10040404",
         967 => x"04040404",
         968 => x"04040410",
         969 => x"10101010",
         970 => x"10104141",
         971 => x"41414141",
         972 => x"01010101",
         973 => x"01010101",
         974 => x"01010101",
         975 => x"01010101",
         976 => x"01010101",
         977 => x"10101010",
         978 => x"10104242",
         979 => x"42424242",
         980 => x"02020202",
         981 => x"02020202",
         982 => x"02020202",
         983 => x"02020202",
         984 => x"02020202",
         985 => x"10101010",
         986 => x"20000000",
         987 => x"00000000",
         988 => x"00000000",
         989 => x"00000000",
         990 => x"00000000",
         991 => x"00000000",
         992 => x"00000000",
         993 => x"00000000",
         994 => x"00000000",
         995 => x"00000000",
         996 => x"00000000",
         997 => x"00000000",
         998 => x"00000000",
         999 => x"00000000",
        1000 => x"00000000",
        1001 => x"00000000",
        1002 => x"00000000",
        1003 => x"00000000",
        1004 => x"00000000",
        1005 => x"00000000",
        1006 => x"00000000",
        1007 => x"00000000",
        1008 => x"00000000",
        1009 => x"00000000",
        1010 => x"00000000",
        1011 => x"00000000",
        1012 => x"00000000",
        1013 => x"00000000",
        1014 => x"00000000",
        1015 => x"00000000",
        1016 => x"00000000",
        1017 => x"00000000",
        1018 => x"00000000"
            );
end package bootrom_image;
