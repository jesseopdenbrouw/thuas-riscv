-- srec2vhdl table generator
-- for input file 'bootloader.srec'
-- date: Fri Sep 27 13:24:06 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package bootrom_image is
    constant bootrom_contents : memory_type := (
           0 => x"97020000",
           1 => x"93820264",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"b7070020",
           9 => x"93870700",
          10 => x"13070500",
          11 => x"3386e740",
          12 => x"63f4e700",
          13 => x"13060000",
          14 => x"93050000",
          15 => x"13050500",
          16 => x"ef004060",
          17 => x"37050020",
          18 => x"b7070020",
          19 => x"93870700",
          20 => x"13070500",
          21 => x"3386e740",
          22 => x"63f4e700",
          23 => x"13060000",
          24 => x"b7150010",
          25 => x"938585f8",
          26 => x"13050500",
          27 => x"ef00405f",
          28 => x"ef009030",
          29 => x"37c50100",
          30 => x"93051000",
          31 => x"13050520",
          32 => x"ef00407e",
          33 => x"ef00902e",
          34 => x"37150010",
          35 => x"130585e2",
          36 => x"ef005002",
          37 => x"732510fc",
          38 => x"37190010",
          39 => x"ef00501d",
          40 => x"130509da",
          41 => x"ef001001",
          42 => x"b70700f0",
          43 => x"1307f03f",
          44 => x"370a1000",
          45 => x"b709a000",
          46 => x"23a2e700",
          47 => x"93041000",
          48 => x"130afaff",
          49 => x"b70a00f0",
          50 => x"93891900",
          51 => x"b3f74401",
          52 => x"639c0700",
          53 => x"1305a002",
          54 => x"ef00c07b",
          55 => x"83a74a00",
          56 => x"93d71700",
          57 => x"23a2fa00",
          58 => x"ef00c05b",
          59 => x"13040500",
          60 => x"63160504",
          61 => x"93841400",
          62 => x"e39a34fd",
          63 => x"b70700f0",
          64 => x"23a20700",
          65 => x"631a0400",
          66 => x"93050000",
          67 => x"13050000",
          68 => x"ef004075",
          69 => x"e7000400",
          70 => x"ef00c059",
          71 => x"1375f50f",
          72 => x"93071002",
          73 => x"6300f502",
          74 => x"93074002",
          75 => x"93040000",
          76 => x"6316f520",
          77 => x"13041000",
          78 => x"6f00c001",
          79 => x"13041000",
          80 => x"6ff0dffb",
          81 => x"37150010",
          82 => x"1305c5e5",
          83 => x"ef008076",
          84 => x"13040000",
          85 => x"93040000",
          86 => x"370a00f0",
          87 => x"130b3005",
          88 => x"930ba004",
          89 => x"130c3002",
          90 => x"93092000",
          91 => x"930ca000",
          92 => x"b71a0010",
          93 => x"83274a00",
          94 => x"93c71700",
          95 => x"2322fa00",
          96 => x"ef004053",
          97 => x"1375f50f",
          98 => x"631e6517",
          99 => x"ef008052",
         100 => x"137df50f",
         101 => x"9307fdfc",
         102 => x"93f7f70f",
         103 => x"63e6f910",
         104 => x"93071003",
         105 => x"631afd04",
         106 => x"13052000",
         107 => x"ef008074",
         108 => x"930dd5ff",
         109 => x"13054000",
         110 => x"ef00c073",
         111 => x"b70601ff",
         112 => x"b705ffff",
         113 => x"130d0500",
         114 => x"b38dad00",
         115 => x"9386f6ff",
         116 => x"9385f50f",
         117 => x"6398ad05",
         118 => x"130da000",
         119 => x"ef00804d",
         120 => x"1375f50f",
         121 => x"e31ca5ff",
         122 => x"e31604f8",
         123 => x"1385cae5",
         124 => x"ef00406c",
         125 => x"6ff01ff8",
         126 => x"93072003",
         127 => x"13052000",
         128 => x"631afd00",
         129 => x"ef00006f",
         130 => x"930dc5ff",
         131 => x"13056000",
         132 => x"6ff09ffa",
         133 => x"ef00006e",
         134 => x"930db5ff",
         135 => x"13058000",
         136 => x"6ff09ff9",
         137 => x"1378cdff",
         138 => x"13052000",
         139 => x"2326b100",
         140 => x"2324d100",
         141 => x"23220101",
         142 => x"ef00c06b",
         143 => x"03284100",
         144 => x"93070500",
         145 => x"37060001",
         146 => x"13753d00",
         147 => x"03270800",
         148 => x"83268100",
         149 => x"8325c100",
         150 => x"93083000",
         151 => x"1306f6ff",
         152 => x"13031000",
         153 => x"63063503",
         154 => x"630a1503",
         155 => x"630c6500",
         156 => x"137707f0",
         157 => x"b3e7e700",
         158 => x"2320f800",
         159 => x"130d1d00",
         160 => x"6ff05ff5",
         161 => x"3377b700",
         162 => x"93978700",
         163 => x"6ff09ffe",
         164 => x"3377d700",
         165 => x"93970701",
         166 => x"6ff0dffd",
         167 => x"3377c700",
         168 => x"93978701",
         169 => x"6ff01ffd",
         170 => x"93079dfc",
         171 => x"93f7f70f",
         172 => x"63e2f904",
         173 => x"13052000",
         174 => x"ef00c063",
         175 => x"93077003",
         176 => x"13058000",
         177 => x"630afd00",
         178 => x"93078003",
         179 => x"13056000",
         180 => x"6304fd00",
         181 => x"13054000",
         182 => x"ef00c061",
         183 => x"93040500",
         184 => x"130da000",
         185 => x"ef00003d",
         186 => x"1375f50f",
         187 => x"e31ca5ff",
         188 => x"6ff09fef",
         189 => x"ef00003c",
         190 => x"1375f50f",
         191 => x"e31c95ff",
         192 => x"6ff09fee",
         193 => x"6310750b",
         194 => x"63180400",
         195 => x"37150010",
         196 => x"1305c5e5",
         197 => x"ef00005a",
         198 => x"93050000",
         199 => x"13050000",
         200 => x"ef004054",
         201 => x"b70700f0",
         202 => x"23a20700",
         203 => x"e7800400",
         204 => x"b70700f0",
         205 => x"1307a00a",
         206 => x"23a2e700",
         207 => x"97020000",
         208 => x"93824223",
         209 => x"73905230",
         210 => x"b7190010",
         211 => x"130509da",
         212 => x"ef004056",
         213 => x"13040000",
         214 => x"371b0010",
         215 => x"b71b0010",
         216 => x"9389d9c9",
         217 => x"b7170010",
         218 => x"138507e6",
         219 => x"ef008054",
         220 => x"93059002",
         221 => x"13054101",
         222 => x"ef00c035",
         223 => x"b7170010",
         224 => x"130a0500",
         225 => x"938547e6",
         226 => x"13054101",
         227 => x"ef00802f",
         228 => x"631e0500",
         229 => x"37150010",
         230 => x"130585e6",
         231 => x"ef008051",
         232 => x"6f00c003",
         233 => x"e31285e5",
         234 => x"6ff09ff8",
         235 => x"b7170010",
         236 => x"938547f5",
         237 => x"13054101",
         238 => x"ef00c02c",
         239 => x"63140502",
         240 => x"93050000",
         241 => x"ef00004a",
         242 => x"b70700f0",
         243 => x"23a20700",
         244 => x"93020000",
         245 => x"73905230",
         246 => x"e7800400",
         247 => x"e3040af8",
         248 => x"6f004018",
         249 => x"b7170010",
         250 => x"13063000",
         251 => x"938587f5",
         252 => x"13054101",
         253 => x"ef001002",
         254 => x"63100504",
         255 => x"93050000",
         256 => x"13057101",
         257 => x"ef00405b",
         258 => x"93773500",
         259 => x"13040500",
         260 => x"63940706",
         261 => x"93058000",
         262 => x"ef00806e",
         263 => x"37150010",
         264 => x"1305c5f5",
         265 => x"ef000049",
         266 => x"03250400",
         267 => x"93058000",
         268 => x"ef00006d",
         269 => x"6ff09ffa",
         270 => x"13063000",
         271 => x"93058bf7",
         272 => x"13054101",
         273 => x"ef00007d",
         274 => x"631e0502",
         275 => x"93050101",
         276 => x"13057101",
         277 => x"ef004056",
         278 => x"93773500",
         279 => x"13040500",
         280 => x"639c0700",
         281 => x"03250101",
         282 => x"93050000",
         283 => x"ef00c054",
         284 => x"2320a400",
         285 => x"6ff09ff6",
         286 => x"37150010",
         287 => x"130505f6",
         288 => x"6ff0dff1",
         289 => x"13063000",
         290 => x"9385cbf7",
         291 => x"13054101",
         292 => x"ef004078",
         293 => x"83474101",
         294 => x"1307e006",
         295 => x"630c0508",
         296 => x"639ae70a",
         297 => x"93773400",
         298 => x"e39807fc",
         299 => x"130c0404",
         300 => x"b71c0010",
         301 => x"371d0010",
         302 => x"930d80ff",
         303 => x"93058000",
         304 => x"13050400",
         305 => x"ef00c063",
         306 => x"1385ccf5",
         307 => x"ef00803e",
         308 => x"83270400",
         309 => x"93058000",
         310 => x"130a8001",
         311 => x"13850700",
         312 => x"2322f100",
         313 => x"ef00c061",
         314 => x"13050df8",
         315 => x"ef00803c",
         316 => x"b70a00ff",
         317 => x"83274100",
         318 => x"33f55701",
         319 => x"33554501",
         320 => x"b3063501",
         321 => x"83c60600",
         322 => x"93f67609",
         323 => x"63800604",
         324 => x"130a8aff",
         325 => x"ef000038",
         326 => x"93da8a00",
         327 => x"e31cbafd",
         328 => x"13044400",
         329 => x"130509da",
         330 => x"ef00c038",
         331 => x"e3188cf8",
         332 => x"6ff05fe3",
         333 => x"e388e7f6",
         334 => x"93050000",
         335 => x"13057101",
         336 => x"ef008047",
         337 => x"13040500",
         338 => x"6ff0dff5",
         339 => x"1305e002",
         340 => x"6ff01ffc",
         341 => x"e3080ae0",
         342 => x"37150010",
         343 => x"130545f8",
         344 => x"ef004035",
         345 => x"130509da",
         346 => x"ef00c034",
         347 => x"6ff09fdf",
         348 => x"130101fb",
         349 => x"23261104",
         350 => x"23245104",
         351 => x"23226104",
         352 => x"23207104",
         353 => x"232e8102",
         354 => x"232c9102",
         355 => x"232aa102",
         356 => x"2328b102",
         357 => x"2326c102",
         358 => x"2324d102",
         359 => x"2322e102",
         360 => x"2320f102",
         361 => x"232e0101",
         362 => x"232c1101",
         363 => x"232ac101",
         364 => x"2328d101",
         365 => x"2326e101",
         366 => x"2324f101",
         367 => x"73241034",
         368 => x"f3242034",
         369 => x"37150010",
         370 => x"130545e1",
         371 => x"ef00802e",
         372 => x"93058000",
         373 => x"13850400",
         374 => x"ef008052",
         375 => x"37150010",
         376 => x"130505da",
         377 => x"ef00002d",
         378 => x"13044400",
         379 => x"73101434",
         380 => x"0324c103",
         381 => x"8320c104",
         382 => x"83228104",
         383 => x"03234104",
         384 => x"83230104",
         385 => x"83248103",
         386 => x"03254103",
         387 => x"83250103",
         388 => x"0326c102",
         389 => x"83268102",
         390 => x"03274102",
         391 => x"83270102",
         392 => x"0328c101",
         393 => x"83288101",
         394 => x"032e4101",
         395 => x"832e0101",
         396 => x"032fc100",
         397 => x"832f8100",
         398 => x"13010105",
         399 => x"73002030",
         400 => x"6f000000",
         401 => x"13030500",
         402 => x"630a0600",
         403 => x"2300b300",
         404 => x"1306f6ff",
         405 => x"13031300",
         406 => x"e31a06fe",
         407 => x"67800000",
         408 => x"13030500",
         409 => x"630e0600",
         410 => x"83830500",
         411 => x"23007300",
         412 => x"1306f6ff",
         413 => x"13031300",
         414 => x"93851500",
         415 => x"e31606fe",
         416 => x"67800000",
         417 => x"03460500",
         418 => x"83c60500",
         419 => x"13051500",
         420 => x"93851500",
         421 => x"6314d600",
         422 => x"e31606fe",
         423 => x"3305d640",
         424 => x"67800000",
         425 => x"b70700f0",
         426 => x"03a54702",
         427 => x"13758500",
         428 => x"67800000",
         429 => x"370700f0",
         430 => x"13070702",
         431 => x"83274700",
         432 => x"93f78700",
         433 => x"e38c07fe",
         434 => x"03258700",
         435 => x"1375f50f",
         436 => x"67800000",
         437 => x"130101fd",
         438 => x"232e3101",
         439 => x"b7190010",
         440 => x"23248102",
         441 => x"23229102",
         442 => x"23202103",
         443 => x"232c4101",
         444 => x"232a5101",
         445 => x"23286101",
         446 => x"23267101",
         447 => x"23261102",
         448 => x"93040500",
         449 => x"13040000",
         450 => x"938909c5",
         451 => x"13095001",
         452 => x"138bf5ff",
         453 => x"130a2000",
         454 => x"930a2001",
         455 => x"b71b0010",
         456 => x"eff05ff9",
         457 => x"1377f50f",
         458 => x"6340e902",
         459 => x"6352ea02",
         460 => x"9307d7ff",
         461 => x"63eefa00",
         462 => x"93972700",
         463 => x"b387f900",
         464 => x"83a70700",
         465 => x"67800700",
         466 => x"9307f007",
         467 => x"630cf706",
         468 => x"6352640f",
         469 => x"9377f50f",
         470 => x"938607fe",
         471 => x"93f6f60f",
         472 => x"1306e005",
         473 => x"e36ed6fa",
         474 => x"b3868400",
         475 => x"2380f600",
         476 => x"13050700",
         477 => x"13041400",
         478 => x"ef00c011",
         479 => x"6ff05ffa",
         480 => x"b3848400",
         481 => x"37150010",
         482 => x"23800400",
         483 => x"130505da",
         484 => x"ef004012",
         485 => x"8320c102",
         486 => x"13050400",
         487 => x"03248102",
         488 => x"83244102",
         489 => x"03290102",
         490 => x"8329c101",
         491 => x"032a8101",
         492 => x"832a4101",
         493 => x"032b0101",
         494 => x"832bc100",
         495 => x"13010103",
         496 => x"67800000",
         497 => x"635a8002",
         498 => x"1305f007",
         499 => x"ef00800c",
         500 => x"1304f4ff",
         501 => x"6ff0dff4",
         502 => x"13854bda",
         503 => x"ef00800d",
         504 => x"eff05fed",
         505 => x"1377f50f",
         506 => x"13040000",
         507 => x"e350e9f4",
         508 => x"9307f007",
         509 => x"e31ef7f4",
         510 => x"23248101",
         511 => x"130c5001",
         512 => x"13057000",
         513 => x"ef000009",
         514 => x"eff0dfea",
         515 => x"1377f50f",
         516 => x"6348ec02",
         517 => x"032c8100",
         518 => x"6ff05ff1",
         519 => x"635a8002",
         520 => x"1305f007",
         521 => x"1304f4ff",
         522 => x"ef00c006",
         523 => x"e31a04fe",
         524 => x"6ff01fef",
         525 => x"13057000",
         526 => x"ef00c005",
         527 => x"6ff05fee",
         528 => x"9307f007",
         529 => x"e30ef7fa",
         530 => x"032c8100",
         531 => x"6ff05ff0",
         532 => x"eff05fe6",
         533 => x"1377f50f",
         534 => x"93075001",
         535 => x"e3d8e7ec",
         536 => x"6ff01ff9",
         537 => x"f32710fc",
         538 => x"63960700",
         539 => x"b7f7fa02",
         540 => x"93870708",
         541 => x"63060500",
         542 => x"33d5a702",
         543 => x"1305f5ff",
         544 => x"b70700f0",
         545 => x"23a6a702",
         546 => x"23a0b702",
         547 => x"23a20702",
         548 => x"67800000",
         549 => x"370700f0",
         550 => x"1375f50f",
         551 => x"13070702",
         552 => x"2324a700",
         553 => x"83274700",
         554 => x"93f70701",
         555 => x"e38c07fe",
         556 => x"67800000",
         557 => x"630e0502",
         558 => x"130101ff",
         559 => x"23248100",
         560 => x"23261100",
         561 => x"13040500",
         562 => x"03450500",
         563 => x"630a0500",
         564 => x"13041400",
         565 => x"eff01ffc",
         566 => x"03450400",
         567 => x"e31a05fe",
         568 => x"8320c100",
         569 => x"03248100",
         570 => x"13010101",
         571 => x"67800000",
         572 => x"67800000",
         573 => x"130101fe",
         574 => x"232e1100",
         575 => x"232c8100",
         576 => x"6350a00a",
         577 => x"23263101",
         578 => x"b7190010",
         579 => x"232a9100",
         580 => x"23282101",
         581 => x"23244101",
         582 => x"13090500",
         583 => x"93040000",
         584 => x"13040000",
         585 => x"9389d9c9",
         586 => x"130a1000",
         587 => x"6f000001",
         588 => x"3364c400",
         589 => x"93841400",
         590 => x"63029904",
         591 => x"eff09fd7",
         592 => x"b387a900",
         593 => x"83c70700",
         594 => x"130605fd",
         595 => x"13144400",
         596 => x"13f74700",
         597 => x"93f64704",
         598 => x"e31c07fc",
         599 => x"93f73700",
         600 => x"e38a06fc",
         601 => x"63944701",
         602 => x"13050502",
         603 => x"130595fa",
         604 => x"93841400",
         605 => x"3364a400",
         606 => x"e31299fc",
         607 => x"8320c101",
         608 => x"13050400",
         609 => x"03248101",
         610 => x"83244101",
         611 => x"03290101",
         612 => x"8329c100",
         613 => x"032a8100",
         614 => x"13010102",
         615 => x"67800000",
         616 => x"13040000",
         617 => x"8320c101",
         618 => x"13050400",
         619 => x"03248101",
         620 => x"13010102",
         621 => x"67800000",
         622 => x"83470500",
         623 => x"37160010",
         624 => x"1306d6c9",
         625 => x"3307f600",
         626 => x"03470700",
         627 => x"93060500",
         628 => x"13758700",
         629 => x"630e0500",
         630 => x"83c71600",
         631 => x"93861600",
         632 => x"3307f600",
         633 => x"03470700",
         634 => x"13758700",
         635 => x"e31605fe",
         636 => x"13754704",
         637 => x"630a0506",
         638 => x"13050000",
         639 => x"13031000",
         640 => x"6f000002",
         641 => x"83c71600",
         642 => x"33e5a800",
         643 => x"93861600",
         644 => x"3307f600",
         645 => x"03470700",
         646 => x"13784704",
         647 => x"63000804",
         648 => x"13784700",
         649 => x"938807fd",
         650 => x"13773700",
         651 => x"13154500",
         652 => x"e31a08fc",
         653 => x"63146700",
         654 => x"93870702",
         655 => x"938797fa",
         656 => x"33e5a700",
         657 => x"83c71600",
         658 => x"93861600",
         659 => x"3307f600",
         660 => x"03470700",
         661 => x"13784704",
         662 => x"e31408fc",
         663 => x"63840500",
         664 => x"23a0d500",
         665 => x"67800000",
         666 => x"13050000",
         667 => x"6ff01fff",
         668 => x"130101fe",
         669 => x"232e1100",
         670 => x"23220100",
         671 => x"23240100",
         672 => x"23260100",
         673 => x"63040506",
         674 => x"232c8100",
         675 => x"93070500",
         676 => x"13040500",
         677 => x"63440504",
         678 => x"13074100",
         679 => x"1306a000",
         680 => x"13089000",
         681 => x"b3f6c702",
         682 => x"13050700",
         683 => x"1307f7ff",
         684 => x"93850700",
         685 => x"93860603",
         686 => x"a305d700",
         687 => x"b3d7c702",
         688 => x"e362b8fe",
         689 => x"3305c500",
         690 => x"eff0dfde",
         691 => x"8320c101",
         692 => x"03248101",
         693 => x"13010102",
         694 => x"67800000",
         695 => x"1305d002",
         696 => x"eff05fdb",
         697 => x"b3078040",
         698 => x"6ff01ffb",
         699 => x"13050003",
         700 => x"eff05fda",
         701 => x"8320c101",
         702 => x"13010102",
         703 => x"67800000",
         704 => x"130101fe",
         705 => x"232e1100",
         706 => x"23220100",
         707 => x"23240100",
         708 => x"23060100",
         709 => x"9387f5ff",
         710 => x"13077000",
         711 => x"6376f700",
         712 => x"93077000",
         713 => x"93058000",
         714 => x"13074100",
         715 => x"b307f700",
         716 => x"b385b740",
         717 => x"13069003",
         718 => x"9376f500",
         719 => x"13870603",
         720 => x"6374e600",
         721 => x"13877605",
         722 => x"2380e700",
         723 => x"9387f7ff",
         724 => x"13554500",
         725 => x"e392f5fe",
         726 => x"13054100",
         727 => x"eff09fd5",
         728 => x"8320c101",
         729 => x"13010102",
         730 => x"67800000",
         731 => x"37150010",
         732 => x"130505db",
         733 => x"6ff01fd4",
         734 => x"130101ff",
         735 => x"23248100",
         736 => x"23229100",
         737 => x"37140010",
         738 => x"b7140010",
         739 => x"938784f8",
         740 => x"130484f8",
         741 => x"3304f440",
         742 => x"23202101",
         743 => x"23261100",
         744 => x"13542440",
         745 => x"938484f8",
         746 => x"13090000",
         747 => x"63108904",
         748 => x"b7140010",
         749 => x"37140010",
         750 => x"938784f8",
         751 => x"130484f8",
         752 => x"3304f440",
         753 => x"13542440",
         754 => x"938484f8",
         755 => x"13090000",
         756 => x"63188902",
         757 => x"8320c100",
         758 => x"03248100",
         759 => x"83244100",
         760 => x"03290100",
         761 => x"13010101",
         762 => x"67800000",
         763 => x"83a70400",
         764 => x"13091900",
         765 => x"93844400",
         766 => x"e7800700",
         767 => x"6ff01ffb",
         768 => x"83a70400",
         769 => x"13091900",
         770 => x"93844400",
         771 => x"e7800700",
         772 => x"6ff01ffc",
         773 => x"630a0602",
         774 => x"1306f6ff",
         775 => x"13070000",
         776 => x"b307e500",
         777 => x"b386e500",
         778 => x"83c70700",
         779 => x"83c60600",
         780 => x"6398d700",
         781 => x"6306c700",
         782 => x"13071700",
         783 => x"e39207fe",
         784 => x"3385d740",
         785 => x"67800000",
         786 => x"13050000",
         787 => x"67800000",
         788 => x"d8070010",
         789 => x"50070010",
         790 => x"50070010",
         791 => x"50070010",
         792 => x"50070010",
         793 => x"c4070010",
         794 => x"50070010",
         795 => x"80070010",
         796 => x"50070010",
         797 => x"50070010",
         798 => x"80070010",
         799 => x"50070010",
         800 => x"50070010",
         801 => x"50070010",
         802 => x"50070010",
         803 => x"50070010",
         804 => x"50070010",
         805 => x"50070010",
         806 => x"1c080010",
         807 => x"00202020",
         808 => x"20202020",
         809 => x"20202828",
         810 => x"28282820",
         811 => x"20202020",
         812 => x"20202020",
         813 => x"20202020",
         814 => x"20202020",
         815 => x"20881010",
         816 => x"10101010",
         817 => x"10101010",
         818 => x"10101010",
         819 => x"10040404",
         820 => x"04040404",
         821 => x"04040410",
         822 => x"10101010",
         823 => x"10104141",
         824 => x"41414141",
         825 => x"01010101",
         826 => x"01010101",
         827 => x"01010101",
         828 => x"01010101",
         829 => x"01010101",
         830 => x"10101010",
         831 => x"10104242",
         832 => x"42424242",
         833 => x"02020202",
         834 => x"02020202",
         835 => x"02020202",
         836 => x"02020202",
         837 => x"02020202",
         838 => x"10101010",
         839 => x"20000000",
         840 => x"00000000",
         841 => x"00000000",
         842 => x"00000000",
         843 => x"00000000",
         844 => x"00000000",
         845 => x"00000000",
         846 => x"00000000",
         847 => x"00000000",
         848 => x"00000000",
         849 => x"00000000",
         850 => x"00000000",
         851 => x"00000000",
         852 => x"00000000",
         853 => x"00000000",
         854 => x"00000000",
         855 => x"00000000",
         856 => x"00000000",
         857 => x"00000000",
         858 => x"00000000",
         859 => x"00000000",
         860 => x"00000000",
         861 => x"00000000",
         862 => x"00000000",
         863 => x"00000000",
         864 => x"00000000",
         865 => x"00000000",
         866 => x"00000000",
         867 => x"00000000",
         868 => x"00000000",
         869 => x"00000000",
         870 => x"00000000",
         871 => x"00000000",
         872 => x"0d0a0000",
         873 => x"3c627265",
         874 => x"616b3e0d",
         875 => x"0a000000",
         876 => x"0d0a5f5f",
         877 => x"5f202020",
         878 => x"20202020",
         879 => x"5f20205f",
         880 => x"5f202020",
         881 => x"205f205c",
         882 => x"202f5f5f",
         883 => x"205f5f20",
         884 => x"0d0a207c",
         885 => x"207c5f7c",
         886 => x"7c207c7c",
         887 => x"5f7c285f",
         888 => x"202d2d2d",
         889 => x"7c5f2920",
         890 => x"56205f5f",
         891 => x"29205f29",
         892 => x"0d0a207c",
         893 => x"207c207c",
         894 => x"7c5f7c7c",
         895 => x"207c5f5f",
         896 => x"29202020",
         897 => x"7c205c20",
         898 => x"20205f5f",
         899 => x"292f5f5f",
         900 => x"0d0a0000",
         901 => x"54726170",
         902 => x"3a206d63",
         903 => x"61757365",
         904 => x"203d2030",
         905 => x"78000000",
         906 => x"0d0a5448",
         907 => x"55415320",
         908 => x"52495343",
         909 => x"2d562042",
         910 => x"6f6f746c",
         911 => x"6f616465",
         912 => x"72207630",
         913 => x"2e362e33",
         914 => x"0d0a436c",
         915 => x"6f636b20",
         916 => x"66726571",
         917 => x"75656e63",
         918 => x"793a2000",
         919 => x"3f0a0000",
         920 => x"3e200000",
         921 => x"68000000",
         922 => x"48656c70",
         923 => x"3a0d0a20",
         924 => x"68202020",
         925 => x"20202020",
         926 => x"20202020",
         927 => x"20202020",
         928 => x"202d2074",
         929 => x"68697320",
         930 => x"68656c70",
         931 => x"0d0a2072",
         932 => x"20202020",
         933 => x"20202020",
         934 => x"20202020",
         935 => x"20202020",
         936 => x"2d207275",
         937 => x"6e206170",
         938 => x"706c6963",
         939 => x"6174696f",
         940 => x"6e0d0a20",
         941 => x"7277203c",
         942 => x"61646472",
         943 => x"3e202020",
         944 => x"20202020",
         945 => x"202d2072",
         946 => x"65616420",
         947 => x"776f7264",
         948 => x"2066726f",
         949 => x"6d206164",
         950 => x"64720d0a",
         951 => x"20777720",
         952 => x"3c616464",
         953 => x"723e203c",
         954 => x"64617461",
         955 => x"3e202d20",
         956 => x"77726974",
         957 => x"6520776f",
         958 => x"72642064",
         959 => x"61746120",
         960 => x"61742061",
         961 => x"6464720d",
         962 => x"0a206477",
         963 => x"203c6164",
         964 => x"64723e20",
         965 => x"20202020",
         966 => x"2020202d",
         967 => x"2064756d",
         968 => x"70203136",
         969 => x"20776f72",
         970 => x"64730d0a",
         971 => x"206e2020",
         972 => x"20202020",
         973 => x"20202020",
         974 => x"20202020",
         975 => x"20202d20",
         976 => x"64756d70",
         977 => x"206e6578",
         978 => x"74203136",
         979 => x"20776f72",
         980 => x"64730000",
         981 => x"72000000",
         982 => x"72772000",
         983 => x"3a200000",
         984 => x"4e6f7420",
         985 => x"6f6e2034",
         986 => x"2d627974",
         987 => x"6520626f",
         988 => x"756e6461",
         989 => x"72792100",
         990 => x"77772000",
         991 => x"64772000",
         992 => x"20200000",
         993 => x"3f3f0000",
         994 => x"00000000"
            );
end package bootrom_image;
