-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Wed Sep  4 12:21:34 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package rom_image is
    constant rom_contents : memory_type := (
           0 => x"97020000",
           1 => x"9382022f",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"13868186",
           8 => x"9387419b",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13858186",
          13 => x"ef104035",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93878186",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"938545e6",
          21 => x"13050500",
          22 => x"ef10c034",
          23 => x"ef10501c",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10c053",
          29 => x"ef10d00f",
          30 => x"6f104048",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef10804c",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"232c4101",
          40 => x"130a0500",
          41 => x"37350000",
          42 => x"130585c7",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"13044100",
          50 => x"ef10404a",
          51 => x"37390000",
          52 => x"9309c1ff",
          53 => x"93070400",
          54 => x"1309c99f",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef10c046",
          65 => x"37350000",
          66 => x"1305c5c8",
          67 => x"ef100046",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef108043",
          78 => x"37350000",
          79 => x"130585c9",
          80 => x"ef10c042",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74708",
          91 => x"b70600f0",
          92 => x"1377f7fe",
          93 => x"23a2e708",
          94 => x"83a74600",
          95 => x"93c71700",
          96 => x"23a2f600",
          97 => x"67800000",
          98 => x"370700f0",
          99 => x"83274700",
         100 => x"93e70720",
         101 => x"2322f700",
         102 => x"6f000000",
         103 => x"b70700f0",
         104 => x"b70500f0",
         105 => x"370500f0",
         106 => x"9387470f",
         107 => x"9385050f",
         108 => x"83a60700",
         109 => x"03a60500",
         110 => x"03a70700",
         111 => x"e31ad7fe",
         112 => x"b7870100",
         113 => x"b70500f0",
         114 => x"1308f0ff",
         115 => x"9387076a",
         116 => x"23ae050f",
         117 => x"b307f600",
         118 => x"b70600f0",
         119 => x"23ac060f",
         120 => x"33b6c700",
         121 => x"23acf60e",
         122 => x"3306e600",
         123 => x"23aec50e",
         124 => x"83274500",
         125 => x"93c72700",
         126 => x"2322f500",
         127 => x"67800000",
         128 => x"b70700f0",
         129 => x"03a74702",
         130 => x"b70600f0",
         131 => x"93870702",
         132 => x"13778700",
         133 => x"630a0700",
         134 => x"03a74600",
         135 => x"13478700",
         136 => x"23a2e600",
         137 => x"83a78700",
         138 => x"67800000",
         139 => x"b70700f0",
         140 => x"03a7470a",
         141 => x"b70600f0",
         142 => x"1377f7f0",
         143 => x"23a2e70a",
         144 => x"83a74600",
         145 => x"93c74700",
         146 => x"23a2f600",
         147 => x"67800000",
         148 => x"b70700f0",
         149 => x"03a74706",
         150 => x"b70600f0",
         151 => x"137777ff",
         152 => x"23a2e706",
         153 => x"83a74600",
         154 => x"93c70701",
         155 => x"23a2f600",
         156 => x"67800000",
         157 => x"b70700f0",
         158 => x"03a74704",
         159 => x"b70600f0",
         160 => x"137777ff",
         161 => x"23a2e704",
         162 => x"83a74600",
         163 => x"93c70702",
         164 => x"23a2f600",
         165 => x"67800000",
         166 => x"b70700f0",
         167 => x"03a74705",
         168 => x"b70600f0",
         169 => x"137777ff",
         170 => x"23aae704",
         171 => x"83a74600",
         172 => x"93c70708",
         173 => x"23a2f600",
         174 => x"67800000",
         175 => x"b70700f0",
         176 => x"23ae0700",
         177 => x"03a74700",
         178 => x"13470704",
         179 => x"23a2e700",
         180 => x"67800000",
         181 => x"370700f0",
         182 => x"b70600f0",
         183 => x"2326070e",
         184 => x"83a74600",
         185 => x"93c70710",
         186 => x"23a2f600",
         187 => x"67800000",
         188 => x"6f000000",
         189 => x"13050000",
         190 => x"67800000",
         191 => x"13050000",
         192 => x"67800000",
         193 => x"130101f7",
         194 => x"23221100",
         195 => x"23242100",
         196 => x"23263100",
         197 => x"23284100",
         198 => x"232a5100",
         199 => x"232c6100",
         200 => x"232e7100",
         201 => x"23208102",
         202 => x"23229102",
         203 => x"2324a102",
         204 => x"2326b102",
         205 => x"2328c102",
         206 => x"232ad102",
         207 => x"232ce102",
         208 => x"232ef102",
         209 => x"23200105",
         210 => x"23221105",
         211 => x"23242105",
         212 => x"23263105",
         213 => x"23284105",
         214 => x"232a5105",
         215 => x"232c6105",
         216 => x"232e7105",
         217 => x"23208107",
         218 => x"23229107",
         219 => x"2324a107",
         220 => x"2326b107",
         221 => x"2328c107",
         222 => x"232ad107",
         223 => x"232ce107",
         224 => x"232ef107",
         225 => x"f3222034",
         226 => x"23205108",
         227 => x"f3221034",
         228 => x"23225108",
         229 => x"83a20200",
         230 => x"23245108",
         231 => x"f3223034",
         232 => x"23265108",
         233 => x"f3272034",
         234 => x"1307b000",
         235 => x"6374f70c",
         236 => x"37070080",
         237 => x"1307d7ff",
         238 => x"b387e700",
         239 => x"13078001",
         240 => x"636ef700",
         241 => x"37370000",
         242 => x"93972700",
         243 => x"130707a1",
         244 => x"b387e700",
         245 => x"83a70700",
         246 => x"67800700",
         247 => x"03258102",
         248 => x"83220108",
         249 => x"63c80200",
         250 => x"f3221034",
         251 => x"93824200",
         252 => x"73901234",
         253 => x"832fc107",
         254 => x"032f8107",
         255 => x"832e4107",
         256 => x"032e0107",
         257 => x"832dc106",
         258 => x"032d8106",
         259 => x"832c4106",
         260 => x"032c0106",
         261 => x"832bc105",
         262 => x"032b8105",
         263 => x"832a4105",
         264 => x"032a0105",
         265 => x"8329c104",
         266 => x"03298104",
         267 => x"83284104",
         268 => x"03280104",
         269 => x"8327c103",
         270 => x"03278103",
         271 => x"83264103",
         272 => x"03260103",
         273 => x"8325c102",
         274 => x"83244102",
         275 => x"03240102",
         276 => x"8323c101",
         277 => x"03238101",
         278 => x"83224101",
         279 => x"03220101",
         280 => x"8321c100",
         281 => x"03218100",
         282 => x"83204100",
         283 => x"13010109",
         284 => x"73002030",
         285 => x"93061000",
         286 => x"e3f2f6f6",
         287 => x"e360f7f6",
         288 => x"37370000",
         289 => x"93972700",
         290 => x"130747a7",
         291 => x"b387e700",
         292 => x"83a70700",
         293 => x"67800700",
         294 => x"eff09fdb",
         295 => x"03258102",
         296 => x"6ff01ff4",
         297 => x"eff01fe3",
         298 => x"03258102",
         299 => x"6ff05ff3",
         300 => x"eff0dfce",
         301 => x"03258102",
         302 => x"6ff09ff2",
         303 => x"eff01fe0",
         304 => x"03258102",
         305 => x"6ff0dff1",
         306 => x"eff0dfc9",
         307 => x"03258102",
         308 => x"6ff01ff1",
         309 => x"eff09fd5",
         310 => x"03258102",
         311 => x"6ff05ff0",
         312 => x"eff01fd2",
         313 => x"03258102",
         314 => x"6ff09fef",
         315 => x"eff0dfda",
         316 => x"03258102",
         317 => x"6ff0dfee",
         318 => x"eff0dfd7",
         319 => x"03258102",
         320 => x"6ff01fee",
         321 => x"13050100",
         322 => x"eff01fb9",
         323 => x"03258102",
         324 => x"6ff01fed",
         325 => x"9307900a",
         326 => x"6380f814",
         327 => x"63d81703",
         328 => x"9307600d",
         329 => x"638ef818",
         330 => x"938808c0",
         331 => x"9307f000",
         332 => x"63e01705",
         333 => x"b7370000",
         334 => x"938747aa",
         335 => x"93982800",
         336 => x"b388f800",
         337 => x"83a70800",
         338 => x"67800700",
         339 => x"938878fc",
         340 => x"93074002",
         341 => x"63ee1701",
         342 => x"b7370000",
         343 => x"938747ae",
         344 => x"93982800",
         345 => x"b388f800",
         346 => x"83a70800",
         347 => x"67800700",
         348 => x"ef10804a",
         349 => x"93078005",
         350 => x"2320f500",
         351 => x"9307f0ff",
         352 => x"13850700",
         353 => x"6ff0dfe5",
         354 => x"b7270000",
         355 => x"23a2f500",
         356 => x"93070000",
         357 => x"13850700",
         358 => x"6ff09fe4",
         359 => x"93070000",
         360 => x"13850700",
         361 => x"6ff0dfe3",
         362 => x"ef100047",
         363 => x"93079000",
         364 => x"2320f500",
         365 => x"9307f0ff",
         366 => x"13850700",
         367 => x"6ff05fe2",
         368 => x"ef108045",
         369 => x"9307f001",
         370 => x"2320f500",
         371 => x"9307f0ff",
         372 => x"13850700",
         373 => x"6ff0dfe0",
         374 => x"ef100044",
         375 => x"9307d000",
         376 => x"2320f500",
         377 => x"9307f0ff",
         378 => x"13850700",
         379 => x"6ff05fdf",
         380 => x"ef108042",
         381 => x"93072000",
         382 => x"2320f500",
         383 => x"9307f0ff",
         384 => x"13850700",
         385 => x"6ff0dfdd",
         386 => x"13090600",
         387 => x"13840500",
         388 => x"635cc000",
         389 => x"b384c500",
         390 => x"eff01fa6",
         391 => x"2300a400",
         392 => x"13041400",
         393 => x"e39a84fe",
         394 => x"13050900",
         395 => x"6ff05fdb",
         396 => x"13090600",
         397 => x"13840500",
         398 => x"e358c0fe",
         399 => x"b384c500",
         400 => x"03450400",
         401 => x"13041400",
         402 => x"eff05fa3",
         403 => x"e39a84fe",
         404 => x"13050900",
         405 => x"6ff0dfd8",
         406 => x"13090000",
         407 => x"93040500",
         408 => x"13040900",
         409 => x"93090900",
         410 => x"93070900",
         411 => x"732410c8",
         412 => x"f32910c0",
         413 => x"f32710c8",
         414 => x"e31af4fe",
         415 => x"37460f00",
         416 => x"13060624",
         417 => x"93060000",
         418 => x"13850900",
         419 => x"93050400",
         420 => x"ef005011",
         421 => x"37460f00",
         422 => x"23a4a400",
         423 => x"13060624",
         424 => x"93060000",
         425 => x"13850900",
         426 => x"93050400",
         427 => x"ef00804c",
         428 => x"23a0a400",
         429 => x"23a2b400",
         430 => x"13050900",
         431 => x"6ff05fd2",
         432 => x"63180500",
         433 => x"1385819b",
         434 => x"13050500",
         435 => x"6ff05fd1",
         436 => x"b7870020",
         437 => x"93870700",
         438 => x"13070040",
         439 => x"b387e740",
         440 => x"e364f5fe",
         441 => x"ef104033",
         442 => x"9307c000",
         443 => x"2320f500",
         444 => x"1305f0ff",
         445 => x"13050500",
         446 => x"6ff09fce",
         447 => x"13030500",
         448 => x"138e0500",
         449 => x"93080000",
         450 => x"63dc0500",
         451 => x"b337a000",
         452 => x"330eb040",
         453 => x"330efe40",
         454 => x"3303a040",
         455 => x"9308f0ff",
         456 => x"63dc0600",
         457 => x"b337c000",
         458 => x"b306d040",
         459 => x"93c8f8ff",
         460 => x"b386f640",
         461 => x"3306c040",
         462 => x"13070600",
         463 => x"13080300",
         464 => x"93070e00",
         465 => x"639c0628",
         466 => x"b7350000",
         467 => x"938585b7",
         468 => x"6376ce0e",
         469 => x"b7060100",
         470 => x"6378d60c",
         471 => x"93360610",
         472 => x"93b61600",
         473 => x"93963600",
         474 => x"3355d600",
         475 => x"b385a500",
         476 => x"83c50500",
         477 => x"13050002",
         478 => x"b386d500",
         479 => x"b305d540",
         480 => x"630cd500",
         481 => x"b317be00",
         482 => x"b356d300",
         483 => x"3317b600",
         484 => x"b3e7f600",
         485 => x"3318b300",
         486 => x"93550701",
         487 => x"33deb702",
         488 => x"13160701",
         489 => x"13560601",
         490 => x"b3f7b702",
         491 => x"13050e00",
         492 => x"3303c603",
         493 => x"93960701",
         494 => x"93570801",
         495 => x"b3e7d700",
         496 => x"63fe6700",
         497 => x"b307f700",
         498 => x"1305feff",
         499 => x"63e8e700",
         500 => x"63f66700",
         501 => x"1305eeff",
         502 => x"b387e700",
         503 => x"b3876740",
         504 => x"33d3b702",
         505 => x"13180801",
         506 => x"13580801",
         507 => x"b3f7b702",
         508 => x"b3066602",
         509 => x"93970701",
         510 => x"3368f800",
         511 => x"93070300",
         512 => x"637cd800",
         513 => x"33080701",
         514 => x"9307f3ff",
         515 => x"6366e800",
         516 => x"6374d800",
         517 => x"9307e3ff",
         518 => x"13150501",
         519 => x"3365f500",
         520 => x"93050000",
         521 => x"6f00000e",
         522 => x"37050001",
         523 => x"93068001",
         524 => x"e37ca6f2",
         525 => x"93060001",
         526 => x"6ff01ff3",
         527 => x"93060000",
         528 => x"630c0600",
         529 => x"b7070100",
         530 => x"637af60c",
         531 => x"93360610",
         532 => x"93b61600",
         533 => x"93963600",
         534 => x"b357d600",
         535 => x"b385f500",
         536 => x"83c70500",
         537 => x"b387d700",
         538 => x"93060002",
         539 => x"b385f640",
         540 => x"6390f60c",
         541 => x"b307ce40",
         542 => x"93051000",
         543 => x"13530701",
         544 => x"b3de6702",
         545 => x"13160701",
         546 => x"13560601",
         547 => x"93560801",
         548 => x"b3f76702",
         549 => x"13850e00",
         550 => x"330ed603",
         551 => x"93970701",
         552 => x"b3e7f600",
         553 => x"63fec701",
         554 => x"b307f700",
         555 => x"1385feff",
         556 => x"63e8e700",
         557 => x"63f6c701",
         558 => x"1385eeff",
         559 => x"b387e700",
         560 => x"b387c741",
         561 => x"33de6702",
         562 => x"13180801",
         563 => x"13580801",
         564 => x"b3f76702",
         565 => x"b306c603",
         566 => x"93970701",
         567 => x"3368f800",
         568 => x"93070e00",
         569 => x"637cd800",
         570 => x"33080701",
         571 => x"9307feff",
         572 => x"6366e800",
         573 => x"6374d800",
         574 => x"9307eeff",
         575 => x"13150501",
         576 => x"3365f500",
         577 => x"638a0800",
         578 => x"b337a000",
         579 => x"b305b040",
         580 => x"b385f540",
         581 => x"3305a040",
         582 => x"67800000",
         583 => x"b7070001",
         584 => x"93068001",
         585 => x"e37af6f2",
         586 => x"93060001",
         587 => x"6ff0dff2",
         588 => x"3317b600",
         589 => x"b356fe00",
         590 => x"13550701",
         591 => x"331ebe00",
         592 => x"b357f300",
         593 => x"b3e7c701",
         594 => x"33dea602",
         595 => x"13160701",
         596 => x"13560601",
         597 => x"3318b300",
         598 => x"b3f6a602",
         599 => x"3303c603",
         600 => x"93950601",
         601 => x"93d60701",
         602 => x"b3e6b600",
         603 => x"93050e00",
         604 => x"63fe6600",
         605 => x"b306d700",
         606 => x"9305feff",
         607 => x"63e8e600",
         608 => x"63f66600",
         609 => x"9305eeff",
         610 => x"b386e600",
         611 => x"b3866640",
         612 => x"33d3a602",
         613 => x"93970701",
         614 => x"93d70701",
         615 => x"b3f6a602",
         616 => x"33066602",
         617 => x"93960601",
         618 => x"b3e7d700",
         619 => x"93060300",
         620 => x"63fec700",
         621 => x"b307f700",
         622 => x"9306f3ff",
         623 => x"63e8e700",
         624 => x"63f6c700",
         625 => x"9306e3ff",
         626 => x"b387e700",
         627 => x"93950501",
         628 => x"b387c740",
         629 => x"b3e5d500",
         630 => x"6ff05fea",
         631 => x"6366de18",
         632 => x"b7070100",
         633 => x"63f4f604",
         634 => x"13b70610",
         635 => x"13371700",
         636 => x"13173700",
         637 => x"b7370000",
         638 => x"b3d5e600",
         639 => x"938787b7",
         640 => x"b387b700",
         641 => x"83c70700",
         642 => x"b387e700",
         643 => x"13070002",
         644 => x"b305f740",
         645 => x"6316f702",
         646 => x"13051000",
         647 => x"e3e4c6ef",
         648 => x"3335c300",
         649 => x"13351500",
         650 => x"6ff0dfed",
         651 => x"b7070001",
         652 => x"13078001",
         653 => x"e3f0f6fc",
         654 => x"13070001",
         655 => x"6ff09ffb",
         656 => x"3357f600",
         657 => x"b396b600",
         658 => x"b366d700",
         659 => x"3357fe00",
         660 => x"331ebe00",
         661 => x"b357f300",
         662 => x"b3e7c701",
         663 => x"13de0601",
         664 => x"335fc703",
         665 => x"13980601",
         666 => x"13580801",
         667 => x"3316b600",
         668 => x"3377c703",
         669 => x"b30ee803",
         670 => x"13150701",
         671 => x"13d70701",
         672 => x"3367a700",
         673 => x"13050f00",
         674 => x"637ed701",
         675 => x"3387e600",
         676 => x"1305ffff",
         677 => x"6368d700",
         678 => x"6376d701",
         679 => x"1305efff",
         680 => x"3307d700",
         681 => x"3307d741",
         682 => x"b35ec703",
         683 => x"93970701",
         684 => x"93d70701",
         685 => x"3377c703",
         686 => x"3308d803",
         687 => x"13170701",
         688 => x"b3e7e700",
         689 => x"13870e00",
         690 => x"63fe0701",
         691 => x"b387f600",
         692 => x"1387feff",
         693 => x"63e8d700",
         694 => x"63f60701",
         695 => x"1387eeff",
         696 => x"b387d700",
         697 => x"13150501",
         698 => x"b70e0100",
         699 => x"3365e500",
         700 => x"9386feff",
         701 => x"3377d500",
         702 => x"b3870741",
         703 => x"b376d600",
         704 => x"13580501",
         705 => x"13560601",
         706 => x"330ed702",
         707 => x"b306d802",
         708 => x"3307c702",
         709 => x"3308c802",
         710 => x"3306d700",
         711 => x"13570e01",
         712 => x"3307c700",
         713 => x"6374d700",
         714 => x"3308d801",
         715 => x"93560701",
         716 => x"b3860601",
         717 => x"63e6d702",
         718 => x"e394d7ce",
         719 => x"b7070100",
         720 => x"9387f7ff",
         721 => x"3377f700",
         722 => x"13170701",
         723 => x"337efe00",
         724 => x"3313b300",
         725 => x"3307c701",
         726 => x"93050000",
         727 => x"e374e3da",
         728 => x"1305f5ff",
         729 => x"6ff0dfcb",
         730 => x"93050000",
         731 => x"13050000",
         732 => x"6ff05fd9",
         733 => x"93080500",
         734 => x"13830500",
         735 => x"13070600",
         736 => x"13080500",
         737 => x"93870500",
         738 => x"63920628",
         739 => x"b7350000",
         740 => x"938585b7",
         741 => x"6376c30e",
         742 => x"b7060100",
         743 => x"6378d60c",
         744 => x"93360610",
         745 => x"93b61600",
         746 => x"93963600",
         747 => x"3355d600",
         748 => x"b385a500",
         749 => x"83c50500",
         750 => x"13050002",
         751 => x"b386d500",
         752 => x"b305d540",
         753 => x"630cd500",
         754 => x"b317b300",
         755 => x"b3d6d800",
         756 => x"3317b600",
         757 => x"b3e7f600",
         758 => x"3398b800",
         759 => x"93550701",
         760 => x"33d3b702",
         761 => x"13160701",
         762 => x"13560601",
         763 => x"b3f7b702",
         764 => x"13050300",
         765 => x"b3086602",
         766 => x"93960701",
         767 => x"93570801",
         768 => x"b3e7d700",
         769 => x"63fe1701",
         770 => x"b307f700",
         771 => x"1305f3ff",
         772 => x"63e8e700",
         773 => x"63f61701",
         774 => x"1305e3ff",
         775 => x"b387e700",
         776 => x"b3871741",
         777 => x"b3d8b702",
         778 => x"13180801",
         779 => x"13580801",
         780 => x"b3f7b702",
         781 => x"b3061603",
         782 => x"93970701",
         783 => x"3368f800",
         784 => x"93870800",
         785 => x"637cd800",
         786 => x"33080701",
         787 => x"9387f8ff",
         788 => x"6366e800",
         789 => x"6374d800",
         790 => x"9387e8ff",
         791 => x"13150501",
         792 => x"3365f500",
         793 => x"93050000",
         794 => x"67800000",
         795 => x"37050001",
         796 => x"93068001",
         797 => x"e37ca6f2",
         798 => x"93060001",
         799 => x"6ff01ff3",
         800 => x"93060000",
         801 => x"630c0600",
         802 => x"b7070100",
         803 => x"6370f60c",
         804 => x"93360610",
         805 => x"93b61600",
         806 => x"93963600",
         807 => x"b357d600",
         808 => x"b385f500",
         809 => x"83c70500",
         810 => x"b387d700",
         811 => x"93060002",
         812 => x"b385f640",
         813 => x"6396f60a",
         814 => x"b307c340",
         815 => x"93051000",
         816 => x"93580701",
         817 => x"33de1703",
         818 => x"13160701",
         819 => x"13560601",
         820 => x"93560801",
         821 => x"b3f71703",
         822 => x"13050e00",
         823 => x"3303c603",
         824 => x"93970701",
         825 => x"b3e7f600",
         826 => x"63fe6700",
         827 => x"b307f700",
         828 => x"1305feff",
         829 => x"63e8e700",
         830 => x"63f66700",
         831 => x"1305eeff",
         832 => x"b387e700",
         833 => x"b3876740",
         834 => x"33d31703",
         835 => x"13180801",
         836 => x"13580801",
         837 => x"b3f71703",
         838 => x"b3066602",
         839 => x"93970701",
         840 => x"3368f800",
         841 => x"93070300",
         842 => x"637cd800",
         843 => x"33080701",
         844 => x"9307f3ff",
         845 => x"6366e800",
         846 => x"6374d800",
         847 => x"9307e3ff",
         848 => x"13150501",
         849 => x"3365f500",
         850 => x"67800000",
         851 => x"b7070001",
         852 => x"93068001",
         853 => x"e374f6f4",
         854 => x"93060001",
         855 => x"6ff01ff4",
         856 => x"3317b600",
         857 => x"b356f300",
         858 => x"13550701",
         859 => x"3313b300",
         860 => x"b3d7f800",
         861 => x"b3e76700",
         862 => x"33d3a602",
         863 => x"13160701",
         864 => x"13560601",
         865 => x"3398b800",
         866 => x"b3f6a602",
         867 => x"b3086602",
         868 => x"93950601",
         869 => x"93d60701",
         870 => x"b3e6b600",
         871 => x"93050300",
         872 => x"63fe1601",
         873 => x"b306d700",
         874 => x"9305f3ff",
         875 => x"63e8e600",
         876 => x"63f61601",
         877 => x"9305e3ff",
         878 => x"b386e600",
         879 => x"b3861641",
         880 => x"b3d8a602",
         881 => x"93970701",
         882 => x"93d70701",
         883 => x"b3f6a602",
         884 => x"33061603",
         885 => x"93960601",
         886 => x"b3e7d700",
         887 => x"93860800",
         888 => x"63fec700",
         889 => x"b307f700",
         890 => x"9386f8ff",
         891 => x"63e8e700",
         892 => x"63f6c700",
         893 => x"9386e8ff",
         894 => x"b387e700",
         895 => x"93950501",
         896 => x"b387c740",
         897 => x"b3e5d500",
         898 => x"6ff09feb",
         899 => x"63e6d518",
         900 => x"b7070100",
         901 => x"63f4f604",
         902 => x"13b70610",
         903 => x"13371700",
         904 => x"13173700",
         905 => x"b7370000",
         906 => x"b3d5e600",
         907 => x"938787b7",
         908 => x"b387b700",
         909 => x"83c70700",
         910 => x"b387e700",
         911 => x"13070002",
         912 => x"b305f740",
         913 => x"6316f702",
         914 => x"13051000",
         915 => x"e3ee66e0",
         916 => x"33b5c800",
         917 => x"13351500",
         918 => x"67800000",
         919 => x"b7070001",
         920 => x"13078001",
         921 => x"e3f0f6fc",
         922 => x"13070001",
         923 => x"6ff09ffb",
         924 => x"3357f600",
         925 => x"b396b600",
         926 => x"b366d700",
         927 => x"3357f300",
         928 => x"3313b300",
         929 => x"b3d7f800",
         930 => x"b3e76700",
         931 => x"13d30601",
         932 => x"b35e6702",
         933 => x"13980601",
         934 => x"13580801",
         935 => x"3316b600",
         936 => x"33776702",
         937 => x"330ed803",
         938 => x"13150701",
         939 => x"13d70701",
         940 => x"3367a700",
         941 => x"13850e00",
         942 => x"637ec701",
         943 => x"3387e600",
         944 => x"1385feff",
         945 => x"6368d700",
         946 => x"6376c701",
         947 => x"1385eeff",
         948 => x"3307d700",
         949 => x"3307c741",
         950 => x"335e6702",
         951 => x"93970701",
         952 => x"93d70701",
         953 => x"33776702",
         954 => x"3308c803",
         955 => x"13170701",
         956 => x"b3e7e700",
         957 => x"13070e00",
         958 => x"63fe0701",
         959 => x"b387f600",
         960 => x"1307feff",
         961 => x"63e8d700",
         962 => x"63f60701",
         963 => x"1307eeff",
         964 => x"b387d700",
         965 => x"13150501",
         966 => x"370e0100",
         967 => x"3365e500",
         968 => x"9306feff",
         969 => x"3377d500",
         970 => x"b3870741",
         971 => x"b376d600",
         972 => x"13580501",
         973 => x"13560601",
         974 => x"3303d702",
         975 => x"b306d802",
         976 => x"3307c702",
         977 => x"3308c802",
         978 => x"3306d700",
         979 => x"13570301",
         980 => x"3307c700",
         981 => x"6374d700",
         982 => x"3308c801",
         983 => x"93560701",
         984 => x"b3860601",
         985 => x"63e6d702",
         986 => x"e39ed7ce",
         987 => x"b7070100",
         988 => x"9387f7ff",
         989 => x"3377f700",
         990 => x"13170701",
         991 => x"3373f300",
         992 => x"b398b800",
         993 => x"33076700",
         994 => x"93050000",
         995 => x"e3fee8cc",
         996 => x"1305f5ff",
         997 => x"6ff01fcd",
         998 => x"93050000",
         999 => x"13050000",
        1000 => x"67800000",
        1001 => x"13080600",
        1002 => x"93070500",
        1003 => x"13870500",
        1004 => x"63960620",
        1005 => x"b7380000",
        1006 => x"938888b7",
        1007 => x"63fcc50c",
        1008 => x"b7060100",
        1009 => x"637ed60a",
        1010 => x"93360610",
        1011 => x"93b61600",
        1012 => x"93963600",
        1013 => x"3353d600",
        1014 => x"b3886800",
        1015 => x"83c80800",
        1016 => x"13030002",
        1017 => x"b386d800",
        1018 => x"b308d340",
        1019 => x"630cd300",
        1020 => x"33971501",
        1021 => x"b356d500",
        1022 => x"33181601",
        1023 => x"33e7e600",
        1024 => x"b3171501",
        1025 => x"13560801",
        1026 => x"b356c702",
        1027 => x"13150801",
        1028 => x"13550501",
        1029 => x"3377c702",
        1030 => x"b386a602",
        1031 => x"93150701",
        1032 => x"13d70701",
        1033 => x"3367b700",
        1034 => x"637ad700",
        1035 => x"3307e800",
        1036 => x"63660701",
        1037 => x"6374d700",
        1038 => x"33070701",
        1039 => x"3307d740",
        1040 => x"b356c702",
        1041 => x"3377c702",
        1042 => x"b386a602",
        1043 => x"93970701",
        1044 => x"13170701",
        1045 => x"93d70701",
        1046 => x"b3e7e700",
        1047 => x"63fad700",
        1048 => x"b307f800",
        1049 => x"63e60701",
        1050 => x"63f4d700",
        1051 => x"b3870701",
        1052 => x"b387d740",
        1053 => x"33d51701",
        1054 => x"93050000",
        1055 => x"67800000",
        1056 => x"37030001",
        1057 => x"93068001",
        1058 => x"e37666f4",
        1059 => x"93060001",
        1060 => x"6ff05ff4",
        1061 => x"93060000",
        1062 => x"630c0600",
        1063 => x"37070100",
        1064 => x"637ee606",
        1065 => x"93360610",
        1066 => x"93b61600",
        1067 => x"93963600",
        1068 => x"3357d600",
        1069 => x"b388e800",
        1070 => x"03c70800",
        1071 => x"3307d700",
        1072 => x"93060002",
        1073 => x"b388e640",
        1074 => x"6394e606",
        1075 => x"3387c540",
        1076 => x"93550801",
        1077 => x"3356b702",
        1078 => x"13150801",
        1079 => x"13550501",
        1080 => x"93d60701",
        1081 => x"3377b702",
        1082 => x"3306a602",
        1083 => x"13170701",
        1084 => x"33e7e600",
        1085 => x"637ac700",
        1086 => x"3307e800",
        1087 => x"63660701",
        1088 => x"6374c700",
        1089 => x"33070701",
        1090 => x"3307c740",
        1091 => x"b356b702",
        1092 => x"3377b702",
        1093 => x"b386a602",
        1094 => x"6ff05ff3",
        1095 => x"37070001",
        1096 => x"93068001",
        1097 => x"e376e6f8",
        1098 => x"93060001",
        1099 => x"6ff05ff8",
        1100 => x"33181601",
        1101 => x"b3d6e500",
        1102 => x"b3171501",
        1103 => x"b3951501",
        1104 => x"3357e500",
        1105 => x"13550801",
        1106 => x"3367b700",
        1107 => x"b3d5a602",
        1108 => x"13130801",
        1109 => x"13530301",
        1110 => x"b3f6a602",
        1111 => x"b3856502",
        1112 => x"13960601",
        1113 => x"93560701",
        1114 => x"b3e6c600",
        1115 => x"63fab600",
        1116 => x"b306d800",
        1117 => x"63e60601",
        1118 => x"63f4b600",
        1119 => x"b3860601",
        1120 => x"b386b640",
        1121 => x"33d6a602",
        1122 => x"13170701",
        1123 => x"13570701",
        1124 => x"b3f6a602",
        1125 => x"33066602",
        1126 => x"93960601",
        1127 => x"3367d700",
        1128 => x"637ac700",
        1129 => x"3307e800",
        1130 => x"63660701",
        1131 => x"6374c700",
        1132 => x"33070701",
        1133 => x"3307c740",
        1134 => x"6ff09ff1",
        1135 => x"63e4d51c",
        1136 => x"37080100",
        1137 => x"63fe0605",
        1138 => x"13b80610",
        1139 => x"13381800",
        1140 => x"13183800",
        1141 => x"b7380000",
        1142 => x"33d30601",
        1143 => x"938888b7",
        1144 => x"b3886800",
        1145 => x"83c80800",
        1146 => x"13030002",
        1147 => x"b3880801",
        1148 => x"33081341",
        1149 => x"63101305",
        1150 => x"63e4b600",
        1151 => x"636cc500",
        1152 => x"3306c540",
        1153 => x"b386d540",
        1154 => x"3337c500",
        1155 => x"93070600",
        1156 => x"3387e640",
        1157 => x"13850700",
        1158 => x"93050700",
        1159 => x"67800000",
        1160 => x"b7080001",
        1161 => x"13088001",
        1162 => x"e3f616fb",
        1163 => x"13080001",
        1164 => x"6ff05ffa",
        1165 => x"b3571601",
        1166 => x"b3960601",
        1167 => x"b3e6d700",
        1168 => x"33d71501",
        1169 => x"13de0601",
        1170 => x"335fc703",
        1171 => x"13930601",
        1172 => x"13530301",
        1173 => x"b3970501",
        1174 => x"b3551501",
        1175 => x"b3e5f500",
        1176 => x"93d70501",
        1177 => x"33160601",
        1178 => x"33150501",
        1179 => x"3377c703",
        1180 => x"b30ee303",
        1181 => x"13170701",
        1182 => x"b3e7e700",
        1183 => x"13070f00",
        1184 => x"63fed701",
        1185 => x"b387f600",
        1186 => x"1307ffff",
        1187 => x"63e8d700",
        1188 => x"63f6d701",
        1189 => x"1307efff",
        1190 => x"b387d700",
        1191 => x"b387d741",
        1192 => x"b3dec703",
        1193 => x"93950501",
        1194 => x"93d50501",
        1195 => x"b3f7c703",
        1196 => x"138e0e00",
        1197 => x"3303d303",
        1198 => x"93970701",
        1199 => x"b3e5f500",
        1200 => x"63fe6500",
        1201 => x"b385b600",
        1202 => x"138efeff",
        1203 => x"63e8d500",
        1204 => x"63f66500",
        1205 => x"138eeeff",
        1206 => x"b385d500",
        1207 => x"93170701",
        1208 => x"370f0100",
        1209 => x"b3e7c701",
        1210 => x"b3856540",
        1211 => x"1303ffff",
        1212 => x"33f76700",
        1213 => x"135e0601",
        1214 => x"93d70701",
        1215 => x"33736600",
        1216 => x"b30e6702",
        1217 => x"33836702",
        1218 => x"3307c703",
        1219 => x"b387c703",
        1220 => x"330e6700",
        1221 => x"13d70e01",
        1222 => x"3307c701",
        1223 => x"63746700",
        1224 => x"b387e701",
        1225 => x"13530701",
        1226 => x"b307f300",
        1227 => x"37030100",
        1228 => x"1303f3ff",
        1229 => x"33776700",
        1230 => x"13170701",
        1231 => x"b3fe6e00",
        1232 => x"3307d701",
        1233 => x"63e6f500",
        1234 => x"639ef500",
        1235 => x"637ce500",
        1236 => x"3306c740",
        1237 => x"3333c700",
        1238 => x"b306d300",
        1239 => x"13070600",
        1240 => x"b387d740",
        1241 => x"3307e540",
        1242 => x"3335e500",
        1243 => x"b385f540",
        1244 => x"b385a540",
        1245 => x"b3981501",
        1246 => x"33570701",
        1247 => x"33e5e800",
        1248 => x"b3d50501",
        1249 => x"67800000",
        1250 => x"13030500",
        1251 => x"630a0600",
        1252 => x"2300b300",
        1253 => x"1306f6ff",
        1254 => x"13031300",
        1255 => x"e31a06fe",
        1256 => x"67800000",
        1257 => x"13030500",
        1258 => x"630e0600",
        1259 => x"83830500",
        1260 => x"23007300",
        1261 => x"1306f6ff",
        1262 => x"13031300",
        1263 => x"93851500",
        1264 => x"e31606fe",
        1265 => x"67800000",
        1266 => x"630c0602",
        1267 => x"13030500",
        1268 => x"93061000",
        1269 => x"636ab500",
        1270 => x"9306f0ff",
        1271 => x"1307f6ff",
        1272 => x"3303e300",
        1273 => x"b385e500",
        1274 => x"83830500",
        1275 => x"23007300",
        1276 => x"1306f6ff",
        1277 => x"3303d300",
        1278 => x"b385d500",
        1279 => x"e31606fe",
        1280 => x"67800000",
        1281 => x"6f000000",
        1282 => x"130101ff",
        1283 => x"23248100",
        1284 => x"13040000",
        1285 => x"23229100",
        1286 => x"23202101",
        1287 => x"23261100",
        1288 => x"93040500",
        1289 => x"13090400",
        1290 => x"93070400",
        1291 => x"732410c8",
        1292 => x"732910c0",
        1293 => x"f32710c8",
        1294 => x"e31af4fe",
        1295 => x"37460f00",
        1296 => x"13060624",
        1297 => x"93060000",
        1298 => x"13050900",
        1299 => x"93050400",
        1300 => x"eff05fb5",
        1301 => x"37460f00",
        1302 => x"23a4a400",
        1303 => x"93050400",
        1304 => x"13050900",
        1305 => x"13060624",
        1306 => x"93060000",
        1307 => x"eff08ff0",
        1308 => x"8320c100",
        1309 => x"03248100",
        1310 => x"23a0a400",
        1311 => x"23a2b400",
        1312 => x"03290100",
        1313 => x"83244100",
        1314 => x"13050000",
        1315 => x"13010101",
        1316 => x"67800000",
        1317 => x"03a78186",
        1318 => x"b7870020",
        1319 => x"93870700",
        1320 => x"93060040",
        1321 => x"b387d740",
        1322 => x"630c0700",
        1323 => x"3305a700",
        1324 => x"63e2a702",
        1325 => x"23a4a186",
        1326 => x"13050700",
        1327 => x"67800000",
        1328 => x"9386819b",
        1329 => x"1387819b",
        1330 => x"23a4d186",
        1331 => x"3305a700",
        1332 => x"e3f2a7fe",
        1333 => x"130101ff",
        1334 => x"23261100",
        1335 => x"ef00c053",
        1336 => x"8320c100",
        1337 => x"9307c000",
        1338 => x"2320f500",
        1339 => x"1307f0ff",
        1340 => x"13050700",
        1341 => x"13010101",
        1342 => x"67800000",
        1343 => x"370700f0",
        1344 => x"13070702",
        1345 => x"83274700",
        1346 => x"93f78700",
        1347 => x"e38c07fe",
        1348 => x"03258700",
        1349 => x"1375f50f",
        1350 => x"67800000",
        1351 => x"f32710fc",
        1352 => x"63960700",
        1353 => x"b7f7fa02",
        1354 => x"93870708",
        1355 => x"63060500",
        1356 => x"33d5a702",
        1357 => x"1305f5ff",
        1358 => x"b70700f0",
        1359 => x"23a6a702",
        1360 => x"23a0b702",
        1361 => x"23a20702",
        1362 => x"67800000",
        1363 => x"370700f0",
        1364 => x"1375f50f",
        1365 => x"13070702",
        1366 => x"2324a700",
        1367 => x"83274700",
        1368 => x"93f70701",
        1369 => x"e38c07fe",
        1370 => x"67800000",
        1371 => x"630e0502",
        1372 => x"130101ff",
        1373 => x"23248100",
        1374 => x"23261100",
        1375 => x"13040500",
        1376 => x"03450500",
        1377 => x"630a0500",
        1378 => x"13041400",
        1379 => x"eff01ffc",
        1380 => x"03450400",
        1381 => x"e31a05fe",
        1382 => x"8320c100",
        1383 => x"03248100",
        1384 => x"13010101",
        1385 => x"67800000",
        1386 => x"67800000",
        1387 => x"130101f8",
        1388 => x"232a9106",
        1389 => x"23282107",
        1390 => x"232e1106",
        1391 => x"232c8106",
        1392 => x"23263107",
        1393 => x"23244107",
        1394 => x"23225107",
        1395 => x"23206107",
        1396 => x"232e7105",
        1397 => x"232c8105",
        1398 => x"232a9105",
        1399 => x"2328a105",
        1400 => x"2326b105",
        1401 => x"13090500",
        1402 => x"93840500",
        1403 => x"f32b00fc",
        1404 => x"b7070008",
        1405 => x"b3fbfb00",
        1406 => x"232c0100",
        1407 => x"232e0100",
        1408 => x"23200102",
        1409 => x"23220102",
        1410 => x"23240102",
        1411 => x"23260102",
        1412 => x"23280102",
        1413 => x"232a0102",
        1414 => x"232c0102",
        1415 => x"232e0102",
        1416 => x"732410fc",
        1417 => x"63160400",
        1418 => x"37f4fa02",
        1419 => x"13040408",
        1420 => x"97f2ffff",
        1421 => x"938242cd",
        1422 => x"73905230",
        1423 => x"37c50100",
        1424 => x"93059000",
        1425 => x"13050520",
        1426 => x"eff05fed",
        1427 => x"b7270000",
        1428 => x"93870771",
        1429 => x"b356f402",
        1430 => x"13561400",
        1431 => x"370700f0",
        1432 => x"1306f6ff",
        1433 => x"b7170300",
        1434 => x"2326c708",
        1435 => x"130e1001",
        1436 => x"938707d4",
        1437 => x"2320c709",
        1438 => x"370600f0",
        1439 => x"37230000",
        1440 => x"1303f370",
        1441 => x"37581200",
        1442 => x"130808f8",
        1443 => x"b70800f0",
        1444 => x"370500f0",
        1445 => x"b70500f0",
        1446 => x"3357f402",
        1447 => x"9387f6ff",
        1448 => x"2328f60a",
        1449 => x"2326660a",
        1450 => x"2320c60b",
        1451 => x"93078070",
        1452 => x"23a0f806",
        1453 => x"b3570403",
        1454 => x"1307f7ff",
        1455 => x"13170701",
        1456 => x"13678700",
        1457 => x"2320e504",
        1458 => x"1307a007",
        1459 => x"9387f7ff",
        1460 => x"93970701",
        1461 => x"93e7c700",
        1462 => x"23a8f504",
        1463 => x"b70700f0",
        1464 => x"23ace700",
        1465 => x"f3224030",
        1466 => x"93e20208",
        1467 => x"73904230",
        1468 => x"f3224030",
        1469 => x"93e28200",
        1470 => x"73904230",
        1471 => x"b7220000",
        1472 => x"93828280",
        1473 => x"73900230",
        1474 => x"b7390000",
        1475 => x"138589c9",
        1476 => x"eff0dfe5",
        1477 => x"1304f9ff",
        1478 => x"63522003",
        1479 => x"1309f0ff",
        1480 => x"03a50400",
        1481 => x"1304f4ff",
        1482 => x"93844400",
        1483 => x"eff01fe4",
        1484 => x"138589c9",
        1485 => x"eff09fe3",
        1486 => x"e31424ff",
        1487 => x"37350000",
        1488 => x"1305c5c9",
        1489 => x"eff09fe2",
        1490 => x"639c0b20",
        1491 => x"37f4eeee",
        1492 => x"b7faeeee",
        1493 => x"b7040010",
        1494 => x"37190000",
        1495 => x"373b0000",
        1496 => x"9384f4ff",
        1497 => x"1304f4ee",
        1498 => x"938aeaee",
        1499 => x"130909e1",
        1500 => x"93090000",
        1501 => x"371c0000",
        1502 => x"130c0c2c",
        1503 => x"130af000",
        1504 => x"6f00c000",
        1505 => x"130cfcff",
        1506 => x"63040c18",
        1507 => x"93050000",
        1508 => x"13058100",
        1509 => x"ef008032",
        1510 => x"e31605fe",
        1511 => x"832c8100",
        1512 => x"8325c100",
        1513 => x"13060900",
        1514 => x"93d7cc01",
        1515 => x"13974500",
        1516 => x"b367f700",
        1517 => x"b3f79700",
        1518 => x"33f79c00",
        1519 => x"13d5f541",
        1520 => x"13d88501",
        1521 => x"3307f700",
        1522 => x"33070701",
        1523 => x"9377d500",
        1524 => x"3307f700",
        1525 => x"33774703",
        1526 => x"937725ff",
        1527 => x"93860900",
        1528 => x"13850c00",
        1529 => x"130cfcff",
        1530 => x"3307f700",
        1531 => x"b387ec40",
        1532 => x"1357f741",
        1533 => x"33b8fc00",
        1534 => x"3387e540",
        1535 => x"33070741",
        1536 => x"b3885703",
        1537 => x"33078702",
        1538 => x"33b88702",
        1539 => x"33071701",
        1540 => x"b3878702",
        1541 => x"33070701",
        1542 => x"1358f741",
        1543 => x"13783800",
        1544 => x"b307f800",
        1545 => x"33b80701",
        1546 => x"3307e800",
        1547 => x"1318e701",
        1548 => x"93d72700",
        1549 => x"b367f800",
        1550 => x"13582740",
        1551 => x"93184800",
        1552 => x"13d3c701",
        1553 => x"33e36800",
        1554 => x"33739300",
        1555 => x"b3f89700",
        1556 => x"135e8801",
        1557 => x"1357f741",
        1558 => x"b3886800",
        1559 => x"b388c801",
        1560 => x"1373d700",
        1561 => x"b3886800",
        1562 => x"b3f84803",
        1563 => x"137727ff",
        1564 => x"139d4700",
        1565 => x"330dfd40",
        1566 => x"131d2d00",
        1567 => x"338dac41",
        1568 => x"b388e800",
        1569 => x"33871741",
        1570 => x"93d8f841",
        1571 => x"33b3e700",
        1572 => x"33081841",
        1573 => x"33086840",
        1574 => x"33088802",
        1575 => x"33035703",
        1576 => x"b3388702",
        1577 => x"33086800",
        1578 => x"33078702",
        1579 => x"33081801",
        1580 => x"9358f841",
        1581 => x"93f83800",
        1582 => x"3387e800",
        1583 => x"b3381701",
        1584 => x"b3880801",
        1585 => x"9398e801",
        1586 => x"13572700",
        1587 => x"33e7e800",
        1588 => x"13184700",
        1589 => x"3307e840",
        1590 => x"13172700",
        1591 => x"b38de740",
        1592 => x"efe0dfe1",
        1593 => x"83260101",
        1594 => x"13070500",
        1595 => x"13080d00",
        1596 => x"93870d00",
        1597 => x"13860c00",
        1598 => x"93054bd0",
        1599 => x"13058101",
        1600 => x"ef00800a",
        1601 => x"13058101",
        1602 => x"eff05fc6",
        1603 => x"e3100ce8",
        1604 => x"63940b00",
        1605 => x"73001000",
        1606 => x"b70700f0",
        1607 => x"9306f00f",
        1608 => x"23a4d706",
        1609 => x"370700f0",
        1610 => x"83260704",
        1611 => x"93050009",
        1612 => x"b70700f0",
        1613 => x"93e60630",
        1614 => x"2320d704",
        1615 => x"2324b704",
        1616 => x"03a60705",
        1617 => x"b70600f0",
        1618 => x"13660630",
        1619 => x"23a8c704",
        1620 => x"23acb704",
        1621 => x"93071000",
        1622 => x"23a6f60e",
        1623 => x"6ff09fe1",
        1624 => x"37350000",
        1625 => x"1305c5cc",
        1626 => x"eff05fc0",
        1627 => x"6ff01fde",
        1628 => x"130101ff",
        1629 => x"23248100",
        1630 => x"23261100",
        1631 => x"93070000",
        1632 => x"13040500",
        1633 => x"63880700",
        1634 => x"93050000",
        1635 => x"97000000",
        1636 => x"e7000000",
        1637 => x"83a7c186",
        1638 => x"63840700",
        1639 => x"e7800700",
        1640 => x"13050400",
        1641 => x"eff01fa6",
        1642 => x"130101f6",
        1643 => x"232af108",
        1644 => x"b7070080",
        1645 => x"9387f7ff",
        1646 => x"232ef100",
        1647 => x"2328f100",
        1648 => x"b707ffff",
        1649 => x"93878720",
        1650 => x"232af100",
        1651 => x"2324a100",
        1652 => x"232ca100",
        1653 => x"03a54186",
        1654 => x"2324c108",
        1655 => x"2326d108",
        1656 => x"13860500",
        1657 => x"93068108",
        1658 => x"93058100",
        1659 => x"232e1106",
        1660 => x"2328e108",
        1661 => x"232c0109",
        1662 => x"232e1109",
        1663 => x"2322d100",
        1664 => x"ef004057",
        1665 => x"83278100",
        1666 => x"23800700",
        1667 => x"8320c107",
        1668 => x"1301010a",
        1669 => x"67800000",
        1670 => x"03a54186",
        1671 => x"67800000",
        1672 => x"130101ff",
        1673 => x"23248100",
        1674 => x"23229100",
        1675 => x"37340000",
        1676 => x"b7340000",
        1677 => x"938744e6",
        1678 => x"130444e6",
        1679 => x"3304f440",
        1680 => x"23202101",
        1681 => x"23261100",
        1682 => x"13542440",
        1683 => x"938444e6",
        1684 => x"13090000",
        1685 => x"63108904",
        1686 => x"b7340000",
        1687 => x"37340000",
        1688 => x"938744e6",
        1689 => x"130444e6",
        1690 => x"3304f440",
        1691 => x"13542440",
        1692 => x"938444e6",
        1693 => x"13090000",
        1694 => x"63188902",
        1695 => x"8320c100",
        1696 => x"03248100",
        1697 => x"83244100",
        1698 => x"03290100",
        1699 => x"13010101",
        1700 => x"67800000",
        1701 => x"83a70400",
        1702 => x"13091900",
        1703 => x"93844400",
        1704 => x"e7800700",
        1705 => x"6ff01ffb",
        1706 => x"83a70400",
        1707 => x"13091900",
        1708 => x"93844400",
        1709 => x"e7800700",
        1710 => x"6ff01ffc",
        1711 => x"13860500",
        1712 => x"93050500",
        1713 => x"03a54186",
        1714 => x"6f00d05a",
        1715 => x"638a050e",
        1716 => x"83a7c5ff",
        1717 => x"130101fe",
        1718 => x"232c8100",
        1719 => x"232e1100",
        1720 => x"1384c5ff",
        1721 => x"63d40700",
        1722 => x"3304f400",
        1723 => x"2326a100",
        1724 => x"ef008031",
        1725 => x"83a78187",
        1726 => x"0325c100",
        1727 => x"639e0700",
        1728 => x"23220400",
        1729 => x"23ac8186",
        1730 => x"03248101",
        1731 => x"8320c101",
        1732 => x"13010102",
        1733 => x"6f00802f",
        1734 => x"6374f402",
        1735 => x"03260400",
        1736 => x"b306c400",
        1737 => x"639ad700",
        1738 => x"83a60700",
        1739 => x"83a74700",
        1740 => x"b386c600",
        1741 => x"2320d400",
        1742 => x"2322f400",
        1743 => x"6ff09ffc",
        1744 => x"13870700",
        1745 => x"83a74700",
        1746 => x"63840700",
        1747 => x"e37af4fe",
        1748 => x"83260700",
        1749 => x"3306d700",
        1750 => x"63188602",
        1751 => x"03260400",
        1752 => x"b386c600",
        1753 => x"2320d700",
        1754 => x"3306d700",
        1755 => x"e39ec7f8",
        1756 => x"03a60700",
        1757 => x"83a74700",
        1758 => x"b306d600",
        1759 => x"2320d700",
        1760 => x"2322f700",
        1761 => x"6ff05ff8",
        1762 => x"6378c400",
        1763 => x"9307c000",
        1764 => x"2320f500",
        1765 => x"6ff05ff7",
        1766 => x"03260400",
        1767 => x"b306c400",
        1768 => x"639ad700",
        1769 => x"83a60700",
        1770 => x"83a74700",
        1771 => x"b386c600",
        1772 => x"2320d400",
        1773 => x"2322f400",
        1774 => x"23228700",
        1775 => x"6ff0dff4",
        1776 => x"67800000",
        1777 => x"130101ff",
        1778 => x"23202101",
        1779 => x"83a74187",
        1780 => x"23248100",
        1781 => x"23229100",
        1782 => x"23261100",
        1783 => x"93040500",
        1784 => x"13840500",
        1785 => x"63980700",
        1786 => x"93050000",
        1787 => x"ef00504d",
        1788 => x"23aaa186",
        1789 => x"93050400",
        1790 => x"13850400",
        1791 => x"ef00504c",
        1792 => x"1309f0ff",
        1793 => x"63122503",
        1794 => x"1304f0ff",
        1795 => x"8320c100",
        1796 => x"13050400",
        1797 => x"03248100",
        1798 => x"83244100",
        1799 => x"03290100",
        1800 => x"13010101",
        1801 => x"67800000",
        1802 => x"13043500",
        1803 => x"1374c4ff",
        1804 => x"e30e85fc",
        1805 => x"b305a440",
        1806 => x"13850400",
        1807 => x"ef005048",
        1808 => x"e31625fd",
        1809 => x"6ff05ffc",
        1810 => x"130101fe",
        1811 => x"232a9100",
        1812 => x"93843500",
        1813 => x"93f4c4ff",
        1814 => x"23282101",
        1815 => x"232e1100",
        1816 => x"232c8100",
        1817 => x"23263101",
        1818 => x"23244101",
        1819 => x"93848400",
        1820 => x"9307c000",
        1821 => x"13090500",
        1822 => x"63f0f40a",
        1823 => x"9304c000",
        1824 => x"63eeb408",
        1825 => x"13050900",
        1826 => x"ef000018",
        1827 => x"83a78187",
        1828 => x"13840700",
        1829 => x"631a040a",
        1830 => x"93850400",
        1831 => x"13050900",
        1832 => x"eff05ff2",
        1833 => x"9307f0ff",
        1834 => x"13040500",
        1835 => x"6316f514",
        1836 => x"03a48187",
        1837 => x"93070400",
        1838 => x"639c0710",
        1839 => x"63040412",
        1840 => x"032a0400",
        1841 => x"93050000",
        1842 => x"13050900",
        1843 => x"330a4401",
        1844 => x"ef00103f",
        1845 => x"6318aa10",
        1846 => x"83270400",
        1847 => x"13050900",
        1848 => x"b384f440",
        1849 => x"93850400",
        1850 => x"eff0dfed",
        1851 => x"9307f0ff",
        1852 => x"630af50e",
        1853 => x"83270400",
        1854 => x"b3879700",
        1855 => x"2320f400",
        1856 => x"83a78187",
        1857 => x"638e070e",
        1858 => x"03a74700",
        1859 => x"6318870c",
        1860 => x"23a20700",
        1861 => x"6f004006",
        1862 => x"e3d404f6",
        1863 => x"9307c000",
        1864 => x"2320f900",
        1865 => x"13050000",
        1866 => x"8320c101",
        1867 => x"03248101",
        1868 => x"83244101",
        1869 => x"03290101",
        1870 => x"8329c100",
        1871 => x"032a8100",
        1872 => x"13010102",
        1873 => x"67800000",
        1874 => x"83260400",
        1875 => x"b3869640",
        1876 => x"63ca0606",
        1877 => x"1307b000",
        1878 => x"637ad704",
        1879 => x"23209400",
        1880 => x"33079400",
        1881 => x"63908704",
        1882 => x"23ace186",
        1883 => x"83274400",
        1884 => x"2320d700",
        1885 => x"2322f700",
        1886 => x"13050900",
        1887 => x"ef000009",
        1888 => x"1305b400",
        1889 => x"93074400",
        1890 => x"137585ff",
        1891 => x"3307f540",
        1892 => x"e30cf5f8",
        1893 => x"3304e400",
        1894 => x"b387a740",
        1895 => x"2320f400",
        1896 => x"6ff09ff8",
        1897 => x"23a2e700",
        1898 => x"6ff05ffc",
        1899 => x"03274400",
        1900 => x"63968700",
        1901 => x"23ace186",
        1902 => x"6ff01ffc",
        1903 => x"23a2e700",
        1904 => x"6ff09ffb",
        1905 => x"93070400",
        1906 => x"03244400",
        1907 => x"6ff09fec",
        1908 => x"13840700",
        1909 => x"83a74700",
        1910 => x"6ff01fee",
        1911 => x"93070700",
        1912 => x"6ff05ff2",
        1913 => x"9307c000",
        1914 => x"2320f900",
        1915 => x"13050900",
        1916 => x"ef00c001",
        1917 => x"6ff01ff3",
        1918 => x"23209500",
        1919 => x"6ff0dff7",
        1920 => x"23220000",
        1921 => x"73001000",
        1922 => x"67800000",
        1923 => x"67800000",
        1924 => x"130101fe",
        1925 => x"23282101",
        1926 => x"03a98500",
        1927 => x"232c8100",
        1928 => x"23263101",
        1929 => x"23225101",
        1930 => x"23206101",
        1931 => x"232e1100",
        1932 => x"232a9100",
        1933 => x"23244101",
        1934 => x"83aa0500",
        1935 => x"13840500",
        1936 => x"130b0600",
        1937 => x"93890600",
        1938 => x"63ec2609",
        1939 => x"8397c500",
        1940 => x"13f70748",
        1941 => x"63040708",
        1942 => x"03274401",
        1943 => x"93043000",
        1944 => x"83a50501",
        1945 => x"b384e402",
        1946 => x"13072000",
        1947 => x"b38aba40",
        1948 => x"130a0500",
        1949 => x"b3c4e402",
        1950 => x"13871600",
        1951 => x"33075701",
        1952 => x"63f4e400",
        1953 => x"93040700",
        1954 => x"93f70740",
        1955 => x"6386070a",
        1956 => x"93850400",
        1957 => x"13050a00",
        1958 => x"eff01fdb",
        1959 => x"13090500",
        1960 => x"630c050a",
        1961 => x"83250401",
        1962 => x"13860a00",
        1963 => x"eff08fcf",
        1964 => x"8357c400",
        1965 => x"93f7f7b7",
        1966 => x"93e70708",
        1967 => x"2316f400",
        1968 => x"23282401",
        1969 => x"232a9400",
        1970 => x"33095901",
        1971 => x"b3845441",
        1972 => x"23202401",
        1973 => x"23249400",
        1974 => x"13890900",
        1975 => x"63f42901",
        1976 => x"13890900",
        1977 => x"03250400",
        1978 => x"13060900",
        1979 => x"93050b00",
        1980 => x"eff08fcd",
        1981 => x"83278400",
        1982 => x"13050000",
        1983 => x"b3872741",
        1984 => x"2324f400",
        1985 => x"83270400",
        1986 => x"b3872701",
        1987 => x"2320f400",
        1988 => x"8320c101",
        1989 => x"03248101",
        1990 => x"83244101",
        1991 => x"03290101",
        1992 => x"8329c100",
        1993 => x"032a8100",
        1994 => x"832a4100",
        1995 => x"032b0100",
        1996 => x"13010102",
        1997 => x"67800000",
        1998 => x"13860400",
        1999 => x"13050a00",
        2000 => x"ef00901c",
        2001 => x"13090500",
        2002 => x"e31c05f6",
        2003 => x"83250401",
        2004 => x"13050a00",
        2005 => x"eff09fb7",
        2006 => x"9307c000",
        2007 => x"2320fa00",
        2008 => x"8357c400",
        2009 => x"1305f0ff",
        2010 => x"93e70704",
        2011 => x"2316f400",
        2012 => x"6ff01ffa",
        2013 => x"83d7c500",
        2014 => x"130101f5",
        2015 => x"2324810a",
        2016 => x"2322910a",
        2017 => x"2320210b",
        2018 => x"232c4109",
        2019 => x"2326110a",
        2020 => x"232e3109",
        2021 => x"232a5109",
        2022 => x"23286109",
        2023 => x"23267109",
        2024 => x"23248109",
        2025 => x"23229109",
        2026 => x"2320a109",
        2027 => x"232eb107",
        2028 => x"93f70708",
        2029 => x"130a0500",
        2030 => x"13890500",
        2031 => x"93040600",
        2032 => x"13840600",
        2033 => x"63880706",
        2034 => x"83a70501",
        2035 => x"63940706",
        2036 => x"93050004",
        2037 => x"eff05fc7",
        2038 => x"2320a900",
        2039 => x"2328a900",
        2040 => x"63160504",
        2041 => x"9307c000",
        2042 => x"2320fa00",
        2043 => x"1305f0ff",
        2044 => x"8320c10a",
        2045 => x"0324810a",
        2046 => x"8324410a",
        2047 => x"0329010a",
        2048 => x"8329c109",
        2049 => x"032a8109",
        2050 => x"832a4109",
        2051 => x"032b0109",
        2052 => x"832bc108",
        2053 => x"032c8108",
        2054 => x"832c4108",
        2055 => x"032d0108",
        2056 => x"832dc107",
        2057 => x"1301010b",
        2058 => x"67800000",
        2059 => x"93070004",
        2060 => x"232af900",
        2061 => x"93070002",
        2062 => x"a304f102",
        2063 => x"93070003",
        2064 => x"23220102",
        2065 => x"2305f102",
        2066 => x"23268100",
        2067 => x"930c5002",
        2068 => x"373b0000",
        2069 => x"b73b0000",
        2070 => x"373d0000",
        2071 => x"372c0000",
        2072 => x"930a0000",
        2073 => x"13840400",
        2074 => x"83470400",
        2075 => x"63840700",
        2076 => x"639c970d",
        2077 => x"b30d9440",
        2078 => x"63069402",
        2079 => x"93860d00",
        2080 => x"13860400",
        2081 => x"93050900",
        2082 => x"13050a00",
        2083 => x"eff05fd8",
        2084 => x"9307f0ff",
        2085 => x"6304f524",
        2086 => x"83274102",
        2087 => x"b387b701",
        2088 => x"2322f102",
        2089 => x"83470400",
        2090 => x"638a0722",
        2091 => x"9307f0ff",
        2092 => x"93041400",
        2093 => x"23280100",
        2094 => x"232e0100",
        2095 => x"232af100",
        2096 => x"232c0100",
        2097 => x"a3090104",
        2098 => x"23240106",
        2099 => x"930d1000",
        2100 => x"83c50400",
        2101 => x"13065000",
        2102 => x"13050bdd",
        2103 => x"ef004077",
        2104 => x"83270101",
        2105 => x"13841400",
        2106 => x"63140506",
        2107 => x"13f70701",
        2108 => x"63060700",
        2109 => x"13070002",
        2110 => x"a309e104",
        2111 => x"13f78700",
        2112 => x"63060700",
        2113 => x"1307b002",
        2114 => x"a309e104",
        2115 => x"83c60400",
        2116 => x"1307a002",
        2117 => x"638ce604",
        2118 => x"8327c101",
        2119 => x"13840400",
        2120 => x"93060000",
        2121 => x"13069000",
        2122 => x"1305a000",
        2123 => x"03470400",
        2124 => x"93051400",
        2125 => x"130707fd",
        2126 => x"637ee608",
        2127 => x"63840604",
        2128 => x"232ef100",
        2129 => x"6f000004",
        2130 => x"13041400",
        2131 => x"6ff0dff1",
        2132 => x"13070bdd",
        2133 => x"3305e540",
        2134 => x"3395ad00",
        2135 => x"b3e7a700",
        2136 => x"2328f100",
        2137 => x"93040400",
        2138 => x"6ff09ff6",
        2139 => x"0327c100",
        2140 => x"93064700",
        2141 => x"03270700",
        2142 => x"2326d100",
        2143 => x"63420704",
        2144 => x"232ee100",
        2145 => x"03470400",
        2146 => x"9307e002",
        2147 => x"6314f708",
        2148 => x"03471400",
        2149 => x"9307a002",
        2150 => x"6318f704",
        2151 => x"8327c100",
        2152 => x"13042400",
        2153 => x"13874700",
        2154 => x"83a70700",
        2155 => x"2326e100",
        2156 => x"63d40700",
        2157 => x"9307f0ff",
        2158 => x"232af100",
        2159 => x"6f008005",
        2160 => x"3307e040",
        2161 => x"93e72700",
        2162 => x"232ee100",
        2163 => x"2328f100",
        2164 => x"6ff05ffb",
        2165 => x"b387a702",
        2166 => x"13840500",
        2167 => x"93061000",
        2168 => x"b387e700",
        2169 => x"6ff09ff4",
        2170 => x"13041400",
        2171 => x"232a0100",
        2172 => x"93060000",
        2173 => x"93070000",
        2174 => x"13069000",
        2175 => x"1305a000",
        2176 => x"03470400",
        2177 => x"93051400",
        2178 => x"130707fd",
        2179 => x"6372e608",
        2180 => x"e39406fa",
        2181 => x"83450400",
        2182 => x"13063000",
        2183 => x"13858bdd",
        2184 => x"ef000063",
        2185 => x"63020502",
        2186 => x"93878bdd",
        2187 => x"3305f540",
        2188 => x"83270101",
        2189 => x"13070004",
        2190 => x"3317a700",
        2191 => x"b3e7e700",
        2192 => x"13041400",
        2193 => x"2328f100",
        2194 => x"83450400",
        2195 => x"13066000",
        2196 => x"1305cddd",
        2197 => x"93041400",
        2198 => x"2304b102",
        2199 => x"ef00405f",
        2200 => x"63080508",
        2201 => x"63980a04",
        2202 => x"03270101",
        2203 => x"8327c100",
        2204 => x"13770710",
        2205 => x"63080702",
        2206 => x"93874700",
        2207 => x"2326f100",
        2208 => x"83274102",
        2209 => x"b3873701",
        2210 => x"2322f102",
        2211 => x"6ff09fdd",
        2212 => x"b387a702",
        2213 => x"13840500",
        2214 => x"93061000",
        2215 => x"b387e700",
        2216 => x"6ff01ff6",
        2217 => x"93877700",
        2218 => x"93f787ff",
        2219 => x"93878700",
        2220 => x"6ff0dffc",
        2221 => x"1307c100",
        2222 => x"93060ce1",
        2223 => x"13060900",
        2224 => x"93050101",
        2225 => x"13050a00",
        2226 => x"97000000",
        2227 => x"e7000000",
        2228 => x"9307f0ff",
        2229 => x"93090500",
        2230 => x"e314f5fa",
        2231 => x"8357c900",
        2232 => x"93f70704",
        2233 => x"e39407d0",
        2234 => x"03254102",
        2235 => x"6ff05fd0",
        2236 => x"1307c100",
        2237 => x"93060ce1",
        2238 => x"13060900",
        2239 => x"93050101",
        2240 => x"13050a00",
        2241 => x"ef00801b",
        2242 => x"6ff09ffc",
        2243 => x"130101fd",
        2244 => x"232a5101",
        2245 => x"83a70501",
        2246 => x"930a0700",
        2247 => x"03a78500",
        2248 => x"23248102",
        2249 => x"23202103",
        2250 => x"232e3101",
        2251 => x"232c4101",
        2252 => x"23261102",
        2253 => x"23229102",
        2254 => x"23286101",
        2255 => x"23267101",
        2256 => x"93090500",
        2257 => x"13840500",
        2258 => x"13090600",
        2259 => x"138a0600",
        2260 => x"63d4e700",
        2261 => x"93070700",
        2262 => x"2320f900",
        2263 => x"03473404",
        2264 => x"63060700",
        2265 => x"93871700",
        2266 => x"2320f900",
        2267 => x"83270400",
        2268 => x"93f70702",
        2269 => x"63880700",
        2270 => x"83270900",
        2271 => x"93872700",
        2272 => x"2320f900",
        2273 => x"83240400",
        2274 => x"93f46400",
        2275 => x"639e0400",
        2276 => x"130b9401",
        2277 => x"930bf0ff",
        2278 => x"8327c400",
        2279 => x"03270900",
        2280 => x"b387e740",
        2281 => x"63c2f408",
        2282 => x"83473404",
        2283 => x"b336f000",
        2284 => x"83270400",
        2285 => x"93f70702",
        2286 => x"6390070c",
        2287 => x"13063404",
        2288 => x"93050a00",
        2289 => x"13850900",
        2290 => x"e7800a00",
        2291 => x"9307f0ff",
        2292 => x"6308f506",
        2293 => x"83270400",
        2294 => x"13074000",
        2295 => x"93040000",
        2296 => x"93f76700",
        2297 => x"639ce700",
        2298 => x"8324c400",
        2299 => x"83270900",
        2300 => x"b384f440",
        2301 => x"63d40400",
        2302 => x"93040000",
        2303 => x"83278400",
        2304 => x"03270401",
        2305 => x"6356f700",
        2306 => x"b387e740",
        2307 => x"b384f400",
        2308 => x"13090000",
        2309 => x"1304a401",
        2310 => x"130bf0ff",
        2311 => x"63902409",
        2312 => x"13050000",
        2313 => x"6f000002",
        2314 => x"93061000",
        2315 => x"13060b00",
        2316 => x"93050a00",
        2317 => x"13850900",
        2318 => x"e7800a00",
        2319 => x"631a7503",
        2320 => x"1305f0ff",
        2321 => x"8320c102",
        2322 => x"03248102",
        2323 => x"83244102",
        2324 => x"03290102",
        2325 => x"8329c101",
        2326 => x"032a8101",
        2327 => x"832a4101",
        2328 => x"032b0101",
        2329 => x"832bc100",
        2330 => x"13010103",
        2331 => x"67800000",
        2332 => x"93841400",
        2333 => x"6ff05ff2",
        2334 => x"3307d400",
        2335 => x"13060003",
        2336 => x"a301c704",
        2337 => x"03475404",
        2338 => x"93871600",
        2339 => x"b307f400",
        2340 => x"93862600",
        2341 => x"a381e704",
        2342 => x"6ff05ff2",
        2343 => x"93061000",
        2344 => x"13060400",
        2345 => x"93050a00",
        2346 => x"13850900",
        2347 => x"e7800a00",
        2348 => x"e30865f9",
        2349 => x"13091900",
        2350 => x"6ff05ff6",
        2351 => x"130101fd",
        2352 => x"23248102",
        2353 => x"23202103",
        2354 => x"232e3101",
        2355 => x"232c4101",
        2356 => x"23261102",
        2357 => x"23229102",
        2358 => x"232a5101",
        2359 => x"23286101",
        2360 => x"138a0600",
        2361 => x"83c68501",
        2362 => x"93078007",
        2363 => x"13090500",
        2364 => x"13840500",
        2365 => x"93090600",
        2366 => x"63eed700",
        2367 => x"93072006",
        2368 => x"13863504",
        2369 => x"63eed700",
        2370 => x"63840628",
        2371 => x"93078005",
        2372 => x"6380f622",
        2373 => x"93042404",
        2374 => x"2301d404",
        2375 => x"6f004004",
        2376 => x"9387d6f9",
        2377 => x"93f7f70f",
        2378 => x"93055001",
        2379 => x"e3e4f5fe",
        2380 => x"b7350000",
        2381 => x"93972700",
        2382 => x"9385c5e0",
        2383 => x"b387b700",
        2384 => x"83a70700",
        2385 => x"67800700",
        2386 => x"83270700",
        2387 => x"93042404",
        2388 => x"93864700",
        2389 => x"83a70700",
        2390 => x"2320d700",
        2391 => x"2301f404",
        2392 => x"93071000",
        2393 => x"6f008026",
        2394 => x"83270400",
        2395 => x"03250700",
        2396 => x"93f60708",
        2397 => x"93054500",
        2398 => x"63860602",
        2399 => x"83270500",
        2400 => x"2320b700",
        2401 => x"37380000",
        2402 => x"63d80700",
        2403 => x"1307d002",
        2404 => x"b307f040",
        2405 => x"a301e404",
        2406 => x"130848de",
        2407 => x"1307a000",
        2408 => x"6f004006",
        2409 => x"93f60704",
        2410 => x"83270500",
        2411 => x"2320b700",
        2412 => x"e38a06fc",
        2413 => x"93970701",
        2414 => x"93d70741",
        2415 => x"6ff09ffc",
        2416 => x"03250400",
        2417 => x"83250700",
        2418 => x"13780508",
        2419 => x"83a70500",
        2420 => x"93854500",
        2421 => x"631a0800",
        2422 => x"13750504",
        2423 => x"63060500",
        2424 => x"93970701",
        2425 => x"93d70701",
        2426 => x"2320b700",
        2427 => x"37380000",
        2428 => x"1307f006",
        2429 => x"130848de",
        2430 => x"639ae614",
        2431 => x"13078000",
        2432 => x"a3010404",
        2433 => x"83264400",
        2434 => x"2324d400",
        2435 => x"63ce0600",
        2436 => x"83250400",
        2437 => x"b3e6d700",
        2438 => x"93040600",
        2439 => x"93f5b5ff",
        2440 => x"2320b400",
        2441 => x"63840602",
        2442 => x"93040600",
        2443 => x"b3f6e702",
        2444 => x"9384f4ff",
        2445 => x"b306d800",
        2446 => x"83c60600",
        2447 => x"2380d400",
        2448 => x"93860700",
        2449 => x"b3d7e702",
        2450 => x"e3f2e6fe",
        2451 => x"93078000",
        2452 => x"6314f702",
        2453 => x"83270400",
        2454 => x"93f71700",
        2455 => x"638e0700",
        2456 => x"03274400",
        2457 => x"83270401",
        2458 => x"63c8e700",
        2459 => x"93070003",
        2460 => x"a38ff4fe",
        2461 => x"9384f4ff",
        2462 => x"33069640",
        2463 => x"2328c400",
        2464 => x"13070a00",
        2465 => x"93860900",
        2466 => x"1306c100",
        2467 => x"93050400",
        2468 => x"13050900",
        2469 => x"eff09fc7",
        2470 => x"930af0ff",
        2471 => x"631e5513",
        2472 => x"1305f0ff",
        2473 => x"8320c102",
        2474 => x"03248102",
        2475 => x"83244102",
        2476 => x"03290102",
        2477 => x"8329c101",
        2478 => x"032a8101",
        2479 => x"832a4101",
        2480 => x"032b0101",
        2481 => x"13010103",
        2482 => x"67800000",
        2483 => x"83270400",
        2484 => x"93e70702",
        2485 => x"2320f400",
        2486 => x"37380000",
        2487 => x"93068007",
        2488 => x"130888df",
        2489 => x"a302d404",
        2490 => x"83260400",
        2491 => x"83250700",
        2492 => x"13f50608",
        2493 => x"83a70500",
        2494 => x"93854500",
        2495 => x"631a0500",
        2496 => x"13f50604",
        2497 => x"63060500",
        2498 => x"93970701",
        2499 => x"93d70701",
        2500 => x"2320b700",
        2501 => x"13f71600",
        2502 => x"63060700",
        2503 => x"93e60602",
        2504 => x"2320d400",
        2505 => x"638c0700",
        2506 => x"13070001",
        2507 => x"6ff05fed",
        2508 => x"37380000",
        2509 => x"130848de",
        2510 => x"6ff0dffa",
        2511 => x"03270400",
        2512 => x"1377f7fd",
        2513 => x"2320e400",
        2514 => x"6ff01ffe",
        2515 => x"1307a000",
        2516 => x"6ff01feb",
        2517 => x"83260400",
        2518 => x"83270700",
        2519 => x"83254401",
        2520 => x"13f80608",
        2521 => x"13854700",
        2522 => x"630a0800",
        2523 => x"2320a700",
        2524 => x"83a70700",
        2525 => x"23a0b700",
        2526 => x"6f008001",
        2527 => x"2320a700",
        2528 => x"93f60604",
        2529 => x"83a70700",
        2530 => x"e38606fe",
        2531 => x"2390b700",
        2532 => x"23280400",
        2533 => x"93040600",
        2534 => x"6ff09fee",
        2535 => x"83270700",
        2536 => x"03264400",
        2537 => x"93050000",
        2538 => x"93864700",
        2539 => x"2320d700",
        2540 => x"83a40700",
        2541 => x"13850400",
        2542 => x"ef008009",
        2543 => x"63060500",
        2544 => x"33059540",
        2545 => x"2322a400",
        2546 => x"83274400",
        2547 => x"2328f400",
        2548 => x"a3010404",
        2549 => x"6ff0dfea",
        2550 => x"83260401",
        2551 => x"13860400",
        2552 => x"93850900",
        2553 => x"13050900",
        2554 => x"e7000a00",
        2555 => x"e30a55eb",
        2556 => x"83270400",
        2557 => x"93f72700",
        2558 => x"63940704",
        2559 => x"8327c100",
        2560 => x"0325c400",
        2561 => x"e350f5ea",
        2562 => x"13850700",
        2563 => x"6ff09fe9",
        2564 => x"93061000",
        2565 => x"13860a00",
        2566 => x"93850900",
        2567 => x"13050900",
        2568 => x"e7000a00",
        2569 => x"e30e65e7",
        2570 => x"93841400",
        2571 => x"8327c400",
        2572 => x"0327c100",
        2573 => x"b387e740",
        2574 => x"e3ccf4fc",
        2575 => x"6ff01ffc",
        2576 => x"93040000",
        2577 => x"930a9401",
        2578 => x"130bf0ff",
        2579 => x"6ff01ffe",
        2580 => x"93f5f50f",
        2581 => x"3306c500",
        2582 => x"6316c500",
        2583 => x"13050000",
        2584 => x"67800000",
        2585 => x"83470500",
        2586 => x"e38cb7fe",
        2587 => x"13051500",
        2588 => x"6ff09ffe",
        2589 => x"130101ff",
        2590 => x"23248100",
        2591 => x"23229100",
        2592 => x"13040500",
        2593 => x"13850500",
        2594 => x"93050600",
        2595 => x"23261100",
        2596 => x"23a80186",
        2597 => x"efe05fb7",
        2598 => x"9307f0ff",
        2599 => x"6318f500",
        2600 => x"83a70187",
        2601 => x"63840700",
        2602 => x"2320f400",
        2603 => x"8320c100",
        2604 => x"03248100",
        2605 => x"83244100",
        2606 => x"13010101",
        2607 => x"67800000",
        2608 => x"130101ff",
        2609 => x"23248100",
        2610 => x"23229100",
        2611 => x"13040500",
        2612 => x"13850500",
        2613 => x"23261100",
        2614 => x"23a80186",
        2615 => x"efe09fbb",
        2616 => x"9307f0ff",
        2617 => x"6318f500",
        2618 => x"83a70187",
        2619 => x"63840700",
        2620 => x"2320f400",
        2621 => x"8320c100",
        2622 => x"03248100",
        2623 => x"83244100",
        2624 => x"13010101",
        2625 => x"67800000",
        2626 => x"130101fe",
        2627 => x"232c8100",
        2628 => x"232e1100",
        2629 => x"232a9100",
        2630 => x"23282101",
        2631 => x"23263101",
        2632 => x"23244101",
        2633 => x"13040600",
        2634 => x"63940502",
        2635 => x"03248101",
        2636 => x"8320c101",
        2637 => x"83244101",
        2638 => x"03290101",
        2639 => x"8329c100",
        2640 => x"032a8100",
        2641 => x"93050600",
        2642 => x"13010102",
        2643 => x"6ff0cfaf",
        2644 => x"63180602",
        2645 => x"eff08f97",
        2646 => x"93040000",
        2647 => x"8320c101",
        2648 => x"03248101",
        2649 => x"03290101",
        2650 => x"8329c100",
        2651 => x"032a8100",
        2652 => x"13850400",
        2653 => x"83244101",
        2654 => x"13010102",
        2655 => x"67800000",
        2656 => x"130a0500",
        2657 => x"93840500",
        2658 => x"ef008005",
        2659 => x"13090500",
        2660 => x"63668500",
        2661 => x"93571500",
        2662 => x"e3e287fc",
        2663 => x"93050400",
        2664 => x"13050a00",
        2665 => x"eff04faa",
        2666 => x"93090500",
        2667 => x"63160500",
        2668 => x"93840900",
        2669 => x"6ff09ffa",
        2670 => x"13060400",
        2671 => x"63748900",
        2672 => x"13060900",
        2673 => x"93850400",
        2674 => x"13850900",
        2675 => x"efe09f9d",
        2676 => x"93850400",
        2677 => x"13050a00",
        2678 => x"eff04f8f",
        2679 => x"6ff05ffd",
        2680 => x"83a7c5ff",
        2681 => x"1385c7ff",
        2682 => x"63d80700",
        2683 => x"b385a500",
        2684 => x"83a70500",
        2685 => x"3305f500",
        2686 => x"67800000",
        2687 => x"30313233",
        2688 => x"34353637",
        2689 => x"38396162",
        2690 => x"63646566",
        2691 => x"00000000",
        2692 => x"a4040000",
        2693 => x"dc030000",
        2694 => x"dc030000",
        2695 => x"dc030000",
        2696 => x"b0040000",
        2697 => x"dc030000",
        2698 => x"dc030000",
        2699 => x"dc030000",
        2700 => x"dc030000",
        2701 => x"dc030000",
        2702 => x"dc030000",
        2703 => x"dc030000",
        2704 => x"dc030000",
        2705 => x"dc030000",
        2706 => x"dc030000",
        2707 => x"bc040000",
        2708 => x"dc030000",
        2709 => x"c8040000",
        2710 => x"d4040000",
        2711 => x"dc030000",
        2712 => x"e0040000",
        2713 => x"ec040000",
        2714 => x"dc030000",
        2715 => x"f8040000",
        2716 => x"98040000",
        2717 => x"dc030000",
        2718 => x"dc030000",
        2719 => x"dc030000",
        2720 => x"04050000",
        2721 => x"dc030000",
        2722 => x"dc030000",
        2723 => x"dc030000",
        2724 => x"dc030000",
        2725 => x"dc030000",
        2726 => x"dc030000",
        2727 => x"dc030000",
        2728 => x"14050000",
        2729 => x"a8050000",
        2730 => x"c0050000",
        2731 => x"f0050000",
        2732 => x"70050000",
        2733 => x"70050000",
        2734 => x"70050000",
        2735 => x"70050000",
        2736 => x"70050000",
        2737 => x"70050000",
        2738 => x"d8050000",
        2739 => x"70050000",
        2740 => x"70050000",
        2741 => x"70050000",
        2742 => x"70050000",
        2743 => x"88050000",
        2744 => x"88050000",
        2745 => x"a8050000",
        2746 => x"70050000",
        2747 => x"70050000",
        2748 => x"70050000",
        2749 => x"70050000",
        2750 => x"9c050000",
        2751 => x"08060000",
        2752 => x"30060000",
        2753 => x"70050000",
        2754 => x"70050000",
        2755 => x"70050000",
        2756 => x"70050000",
        2757 => x"70050000",
        2758 => x"70050000",
        2759 => x"70050000",
        2760 => x"70050000",
        2761 => x"70050000",
        2762 => x"70050000",
        2763 => x"70050000",
        2764 => x"70050000",
        2765 => x"70050000",
        2766 => x"70050000",
        2767 => x"88050000",
        2768 => x"88050000",
        2769 => x"70050000",
        2770 => x"70050000",
        2771 => x"70050000",
        2772 => x"70050000",
        2773 => x"70050000",
        2774 => x"70050000",
        2775 => x"70050000",
        2776 => x"70050000",
        2777 => x"70050000",
        2778 => x"70050000",
        2779 => x"70050000",
        2780 => x"70050000",
        2781 => x"9c050000",
        2782 => x"00010202",
        2783 => x"03030303",
        2784 => x"04040404",
        2785 => x"04040404",
        2786 => x"05050505",
        2787 => x"05050505",
        2788 => x"05050505",
        2789 => x"05050505",
        2790 => x"06060606",
        2791 => x"06060606",
        2792 => x"06060606",
        2793 => x"06060606",
        2794 => x"06060606",
        2795 => x"06060606",
        2796 => x"06060606",
        2797 => x"06060606",
        2798 => x"07070707",
        2799 => x"07070707",
        2800 => x"07070707",
        2801 => x"07070707",
        2802 => x"07070707",
        2803 => x"07070707",
        2804 => x"07070707",
        2805 => x"07070707",
        2806 => x"07070707",
        2807 => x"07070707",
        2808 => x"07070707",
        2809 => x"07070707",
        2810 => x"07070707",
        2811 => x"07070707",
        2812 => x"07070707",
        2813 => x"07070707",
        2814 => x"08080808",
        2815 => x"08080808",
        2816 => x"08080808",
        2817 => x"08080808",
        2818 => x"08080808",
        2819 => x"08080808",
        2820 => x"08080808",
        2821 => x"08080808",
        2822 => x"08080808",
        2823 => x"08080808",
        2824 => x"08080808",
        2825 => x"08080808",
        2826 => x"08080808",
        2827 => x"08080808",
        2828 => x"08080808",
        2829 => x"08080808",
        2830 => x"08080808",
        2831 => x"08080808",
        2832 => x"08080808",
        2833 => x"08080808",
        2834 => x"08080808",
        2835 => x"08080808",
        2836 => x"08080808",
        2837 => x"08080808",
        2838 => x"08080808",
        2839 => x"08080808",
        2840 => x"08080808",
        2841 => x"08080808",
        2842 => x"08080808",
        2843 => x"08080808",
        2844 => x"08080808",
        2845 => x"08080808",
        2846 => x"0d0a4542",
        2847 => x"5245414b",
        2848 => x"21206d65",
        2849 => x"7063203d",
        2850 => x"20000000",
        2851 => x"20696e73",
        2852 => x"6e203d20",
        2853 => x"00000000",
        2854 => x"0d0a0000",
        2855 => x"0d0a0a44",
        2856 => x"6973706c",
        2857 => x"6179696e",
        2858 => x"67207468",
        2859 => x"65207469",
        2860 => x"6d652070",
        2861 => x"61737365",
        2862 => x"64207369",
        2863 => x"6e636520",
        2864 => x"72657365",
        2865 => x"740d0a0a",
        2866 => x"00000000",
        2867 => x"4f6e2d63",
        2868 => x"68697020",
        2869 => x"64656275",
        2870 => x"67676572",
        2871 => x"20666f75",
        2872 => x"6e642c20",
        2873 => x"736b6970",
        2874 => x"70696e67",
        2875 => x"20454252",
        2876 => x"45414b20",
        2877 => x"696e7374",
        2878 => x"72756374",
        2879 => x"696f6e0d",
        2880 => x"0a0d0a00",
        2881 => x"2530356c",
        2882 => x"643a2530",
        2883 => x"366c6420",
        2884 => x"20202530",
        2885 => x"326c643a",
        2886 => x"2530326c",
        2887 => x"643a2530",
        2888 => x"326c640d",
        2889 => x"00000000",
        2890 => x"696e7465",
        2891 => x"72727570",
        2892 => x"745f6469",
        2893 => x"72656374",
        2894 => x"00000000",
        2895 => x"54485541",
        2896 => x"53205249",
        2897 => x"53432d56",
        2898 => x"20525633",
        2899 => x"32494d20",
        2900 => x"62617265",
        2901 => x"206d6574",
        2902 => x"616c2070",
        2903 => x"726f6365",
        2904 => x"73736f72",
        2905 => x"00000000",
        2906 => x"54686520",
        2907 => x"48616775",
        2908 => x"6520556e",
        2909 => x"69766572",
        2910 => x"73697479",
        2911 => x"206f6620",
        2912 => x"4170706c",
        2913 => x"69656420",
        2914 => x"53636965",
        2915 => x"6e636573",
        2916 => x"00000000",
        2917 => x"44657061",
        2918 => x"72746d65",
        2919 => x"6e74206f",
        2920 => x"6620456c",
        2921 => x"65637472",
        2922 => x"6963616c",
        2923 => x"20456e67",
        2924 => x"696e6565",
        2925 => x"72696e67",
        2926 => x"00000000",
        2927 => x"4a2e452e",
        2928 => x"4a2e206f",
        2929 => x"70206465",
        2930 => x"6e204272",
        2931 => x"6f757700",
        2932 => x"232d302b",
        2933 => x"20000000",
        2934 => x"686c4c00",
        2935 => x"65666745",
        2936 => x"46470000",
        2937 => x"30313233",
        2938 => x"34353637",
        2939 => x"38394142",
        2940 => x"43444546",
        2941 => x"00000000",
        2942 => x"30313233",
        2943 => x"34353637",
        2944 => x"38396162",
        2945 => x"63646566",
        2946 => x"00000000",
        2947 => x"48250000",
        2948 => x"68250000",
        2949 => x"14250000",
        2950 => x"14250000",
        2951 => x"14250000",
        2952 => x"14250000",
        2953 => x"68250000",
        2954 => x"14250000",
        2955 => x"14250000",
        2956 => x"14250000",
        2957 => x"14250000",
        2958 => x"54270000",
        2959 => x"c0250000",
        2960 => x"cc260000",
        2961 => x"14250000",
        2962 => x"14250000",
        2963 => x"9c270000",
        2964 => x"14250000",
        2965 => x"c0250000",
        2966 => x"14250000",
        2967 => x"14250000",
        2968 => x"d8260000",
        2969 => x"282d0000",
        2970 => x"3c2d0000",
        2971 => x"682d0000",
        2972 => x"942d0000",
        2973 => x"bc2d0000",
        2974 => x"00000000",
        2975 => x"00000000",
        2976 => x"7c000020",
        2977 => x"e4000020",
        2978 => x"4c010020",
        2979 => x"00000000",
        2980 => x"00000000",
        2981 => x"00000000",
        2982 => x"00000000",
        2983 => x"00000000",
        2984 => x"00000000",
        2985 => x"00000000",
        2986 => x"00000000",
        2987 => x"00000000",
        2988 => x"00000000",
        2989 => x"00000000",
        2990 => x"00000000",
        2991 => x"00000000",
        2992 => x"00000000",
        2993 => x"00000000",
        2994 => x"18000020",
        2995 => x"00000000"
            );
end package rom_image;
