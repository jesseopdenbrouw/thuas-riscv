-- srec2vhdl table generator
-- for input file 'bootloader.srec'
-- date: Mon Apr  1 13:08:27 2024


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package bootrom_image is
    constant bootrom_contents : memory_type := (
           0 => x"97020000",
           1 => x"93820264",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"37050020",
           8 => x"b7070020",
           9 => x"93870700",
          10 => x"13070500",
          11 => x"3386e740",
          12 => x"63f4e700",
          13 => x"13060000",
          14 => x"93050000",
          15 => x"13050500",
          16 => x"ef004060",
          17 => x"37050020",
          18 => x"b7070020",
          19 => x"93870700",
          20 => x"13070500",
          21 => x"3386e740",
          22 => x"63f4e700",
          23 => x"13060000",
          24 => x"b7150010",
          25 => x"938585f1",
          26 => x"13050500",
          27 => x"ef00405f",
          28 => x"ef00902f",
          29 => x"37c50100",
          30 => x"93051000",
          31 => x"13050520",
          32 => x"ef00407e",
          33 => x"37150010",
          34 => x"130545db",
          35 => x"ef005002",
          36 => x"37150010",
          37 => x"130585dd",
          38 => x"ef009001",
          39 => x"732510fc",
          40 => x"37190010",
          41 => x"ef00901c",
          42 => x"130509d9",
          43 => x"ef005000",
          44 => x"b70700f0",
          45 => x"1307f03f",
          46 => x"370a1000",
          47 => x"b709a000",
          48 => x"23a2e700",
          49 => x"93041000",
          50 => x"130afaff",
          51 => x"b70a00f0",
          52 => x"93891900",
          53 => x"b3f74401",
          54 => x"639c0700",
          55 => x"1305a002",
          56 => x"ef00007b",
          57 => x"83a74a00",
          58 => x"93d71700",
          59 => x"23a2fa00",
          60 => x"ef00405b",
          61 => x"13040500",
          62 => x"63160504",
          63 => x"93841400",
          64 => x"e39a34fd",
          65 => x"b70700f0",
          66 => x"23a20700",
          67 => x"631a0400",
          68 => x"93050000",
          69 => x"13050000",
          70 => x"ef00c074",
          71 => x"e7000400",
          72 => x"ef004059",
          73 => x"1375f50f",
          74 => x"93071002",
          75 => x"6300f502",
          76 => x"93074002",
          77 => x"93040000",
          78 => x"6316f520",
          79 => x"13041000",
          80 => x"6f00c001",
          81 => x"13041000",
          82 => x"6ff0dffb",
          83 => x"37150010",
          84 => x"1305c5de",
          85 => x"ef00c075",
          86 => x"13040000",
          87 => x"93040000",
          88 => x"370a00f0",
          89 => x"130b3005",
          90 => x"930ba004",
          91 => x"130c3002",
          92 => x"93092000",
          93 => x"930ca000",
          94 => x"b71a0010",
          95 => x"83274a00",
          96 => x"93c71700",
          97 => x"2322fa00",
          98 => x"ef00c052",
          99 => x"1375f50f",
         100 => x"631e6517",
         101 => x"ef000052",
         102 => x"137df50f",
         103 => x"9307fdfc",
         104 => x"93f7f70f",
         105 => x"63e6f910",
         106 => x"93071003",
         107 => x"631afd04",
         108 => x"13052000",
         109 => x"ef00c073",
         110 => x"930dd5ff",
         111 => x"13054000",
         112 => x"ef000073",
         113 => x"b70601ff",
         114 => x"b705ffff",
         115 => x"130d0500",
         116 => x"b38dad00",
         117 => x"9386f6ff",
         118 => x"9385f50f",
         119 => x"6398ad05",
         120 => x"130da000",
         121 => x"ef00004d",
         122 => x"1375f50f",
         123 => x"e31ca5ff",
         124 => x"e31604f8",
         125 => x"1385cade",
         126 => x"ef00806b",
         127 => x"6ff01ff8",
         128 => x"93072003",
         129 => x"13052000",
         130 => x"631afd00",
         131 => x"ef00406e",
         132 => x"930dc5ff",
         133 => x"13056000",
         134 => x"6ff09ffa",
         135 => x"ef00406d",
         136 => x"930db5ff",
         137 => x"13058000",
         138 => x"6ff09ff9",
         139 => x"1378cdff",
         140 => x"13052000",
         141 => x"2326b100",
         142 => x"2324d100",
         143 => x"23220101",
         144 => x"ef00006b",
         145 => x"03284100",
         146 => x"93070500",
         147 => x"37060001",
         148 => x"13753d00",
         149 => x"03270800",
         150 => x"83268100",
         151 => x"8325c100",
         152 => x"93083000",
         153 => x"1306f6ff",
         154 => x"13031000",
         155 => x"63063503",
         156 => x"630a1503",
         157 => x"630c6500",
         158 => x"137707f0",
         159 => x"b3e7e700",
         160 => x"2320f800",
         161 => x"130d1d00",
         162 => x"6ff05ff5",
         163 => x"3377b700",
         164 => x"93978700",
         165 => x"6ff09ffe",
         166 => x"3377d700",
         167 => x"93970701",
         168 => x"6ff0dffd",
         169 => x"3377c700",
         170 => x"93978701",
         171 => x"6ff01ffd",
         172 => x"93079dfc",
         173 => x"93f7f70f",
         174 => x"63e2f904",
         175 => x"13052000",
         176 => x"ef000063",
         177 => x"93077003",
         178 => x"13058000",
         179 => x"630afd00",
         180 => x"93078003",
         181 => x"13056000",
         182 => x"6304fd00",
         183 => x"13054000",
         184 => x"ef000061",
         185 => x"93040500",
         186 => x"130da000",
         187 => x"ef00803c",
         188 => x"1375f50f",
         189 => x"e31ca5ff",
         190 => x"6ff09fef",
         191 => x"ef00803b",
         192 => x"1375f50f",
         193 => x"e31c95ff",
         194 => x"6ff09fee",
         195 => x"631e7509",
         196 => x"63180400",
         197 => x"37150010",
         198 => x"1305c5de",
         199 => x"ef004059",
         200 => x"93050000",
         201 => x"13050000",
         202 => x"ef00c053",
         203 => x"b70700f0",
         204 => x"23a20700",
         205 => x"e7800400",
         206 => x"b70700f0",
         207 => x"1307a00a",
         208 => x"23a2e700",
         209 => x"97020000",
         210 => x"9382c222",
         211 => x"73905230",
         212 => x"b7190010",
         213 => x"130509d9",
         214 => x"ef008055",
         215 => x"13040000",
         216 => x"b71b0010",
         217 => x"9389d9c8",
         218 => x"b7170010",
         219 => x"138507df",
         220 => x"ef000054",
         221 => x"93059002",
         222 => x"13054101",
         223 => x"ef008035",
         224 => x"b7170010",
         225 => x"130a0500",
         226 => x"938547df",
         227 => x"13054101",
         228 => x"ef00402f",
         229 => x"631e0500",
         230 => x"37150010",
         231 => x"130585df",
         232 => x"ef000051",
         233 => x"6f00c003",
         234 => x"e31485e5",
         235 => x"6ff0dff8",
         236 => x"b7170010",
         237 => x"938547ee",
         238 => x"13054101",
         239 => x"ef00802c",
         240 => x"63140502",
         241 => x"93050000",
         242 => x"ef00c049",
         243 => x"b70700f0",
         244 => x"23a20700",
         245 => x"93020000",
         246 => x"73905230",
         247 => x"e7800400",
         248 => x"e3040af8",
         249 => x"6f000018",
         250 => x"b7170010",
         251 => x"13063000",
         252 => x"938587ee",
         253 => x"13054101",
         254 => x"ef00d000",
         255 => x"63100504",
         256 => x"93050000",
         257 => x"13057101",
         258 => x"ef00c05a",
         259 => x"93773500",
         260 => x"13040500",
         261 => x"63960706",
         262 => x"93058000",
         263 => x"ef00006e",
         264 => x"37150010",
         265 => x"1305c5ee",
         266 => x"ef008048",
         267 => x"03250400",
         268 => x"93058000",
         269 => x"ef00806c",
         270 => x"6ff09ffa",
         271 => x"b7170010",
         272 => x"13063000",
         273 => x"938587f0",
         274 => x"13054101",
         275 => x"ef00807b",
         276 => x"631e0502",
         277 => x"93050101",
         278 => x"13057101",
         279 => x"ef008055",
         280 => x"93773500",
         281 => x"13040500",
         282 => x"639c0700",
         283 => x"03250101",
         284 => x"93050000",
         285 => x"ef000054",
         286 => x"2320a400",
         287 => x"6ff05ff6",
         288 => x"37150010",
         289 => x"130505ef",
         290 => x"6ff09ff1",
         291 => x"13063000",
         292 => x"9385cbf0",
         293 => x"13054101",
         294 => x"ef00c076",
         295 => x"83474101",
         296 => x"1307e006",
         297 => x"63080508",
         298 => x"6396e70a",
         299 => x"93773400",
         300 => x"e39807fc",
         301 => x"130c0404",
         302 => x"b71c0010",
         303 => x"371d0010",
         304 => x"930d80ff",
         305 => x"93058000",
         306 => x"13050400",
         307 => x"ef000063",
         308 => x"1385ccee",
         309 => x"ef00c03d",
         310 => x"032a0400",
         311 => x"93058000",
         312 => x"930a8001",
         313 => x"13050a00",
         314 => x"ef004061",
         315 => x"13050df1",
         316 => x"ef00003c",
         317 => x"370b00ff",
         318 => x"33756a01",
         319 => x"33555501",
         320 => x"b3063501",
         321 => x"83c60600",
         322 => x"93f67609",
         323 => x"63800604",
         324 => x"938a8aff",
         325 => x"ef00c037",
         326 => x"135b8b00",
         327 => x"e39ebafd",
         328 => x"13044400",
         329 => x"130509d9",
         330 => x"ef008038",
         331 => x"e31c8cf8",
         332 => x"6ff09fe3",
         333 => x"e38ce7f6",
         334 => x"93050000",
         335 => x"13057101",
         336 => x"ef004047",
         337 => x"13040500",
         338 => x"6ff05ff6",
         339 => x"1305e002",
         340 => x"6ff01ffc",
         341 => x"e30a0ae0",
         342 => x"37150010",
         343 => x"130545f1",
         344 => x"ef000035",
         345 => x"130509d9",
         346 => x"ef008034",
         347 => x"6ff0dfdf",
         348 => x"130101fb",
         349 => x"23261104",
         350 => x"23245104",
         351 => x"23226104",
         352 => x"23207104",
         353 => x"232e8102",
         354 => x"232c9102",
         355 => x"232aa102",
         356 => x"2328b102",
         357 => x"2326c102",
         358 => x"2324d102",
         359 => x"2322e102",
         360 => x"2320f102",
         361 => x"232e0101",
         362 => x"232c1101",
         363 => x"232ac101",
         364 => x"2328d101",
         365 => x"2326e101",
         366 => x"2324f101",
         367 => x"73241034",
         368 => x"f3242034",
         369 => x"37150010",
         370 => x"130505da",
         371 => x"ef00402e",
         372 => x"93058000",
         373 => x"13850400",
         374 => x"ef004052",
         375 => x"37150010",
         376 => x"130505d9",
         377 => x"ef00c02c",
         378 => x"13044400",
         379 => x"73101434",
         380 => x"0324c103",
         381 => x"8320c104",
         382 => x"83228104",
         383 => x"03234104",
         384 => x"83230104",
         385 => x"83248103",
         386 => x"03254103",
         387 => x"83250103",
         388 => x"0326c102",
         389 => x"83268102",
         390 => x"03274102",
         391 => x"83270102",
         392 => x"0328c101",
         393 => x"83288101",
         394 => x"032e4101",
         395 => x"832e0101",
         396 => x"032fc100",
         397 => x"832f8100",
         398 => x"13010105",
         399 => x"73002030",
         400 => x"6f000000",
         401 => x"13030500",
         402 => x"630a0600",
         403 => x"2300b300",
         404 => x"1306f6ff",
         405 => x"13031300",
         406 => x"e31a06fe",
         407 => x"67800000",
         408 => x"13030500",
         409 => x"630e0600",
         410 => x"83830500",
         411 => x"23007300",
         412 => x"1306f6ff",
         413 => x"13031300",
         414 => x"93851500",
         415 => x"e31606fe",
         416 => x"67800000",
         417 => x"03460500",
         418 => x"83c60500",
         419 => x"13051500",
         420 => x"93851500",
         421 => x"6314d600",
         422 => x"e31606fe",
         423 => x"3305d640",
         424 => x"67800000",
         425 => x"b70700f0",
         426 => x"03a54702",
         427 => x"13758500",
         428 => x"67800000",
         429 => x"370700f0",
         430 => x"13070702",
         431 => x"83274700",
         432 => x"93f78700",
         433 => x"e38c07fe",
         434 => x"03258700",
         435 => x"1375f50f",
         436 => x"67800000",
         437 => x"130101fd",
         438 => x"232e3101",
         439 => x"b7190010",
         440 => x"23248102",
         441 => x"23229102",
         442 => x"23202103",
         443 => x"232c4101",
         444 => x"232a5101",
         445 => x"23286101",
         446 => x"23267101",
         447 => x"23261102",
         448 => x"93040500",
         449 => x"13040000",
         450 => x"938909c4",
         451 => x"13095001",
         452 => x"138bf5ff",
         453 => x"130a2000",
         454 => x"930a2001",
         455 => x"b71b0010",
         456 => x"eff05ff9",
         457 => x"1377f50f",
         458 => x"6340e902",
         459 => x"6352ea02",
         460 => x"9307d7ff",
         461 => x"63eefa00",
         462 => x"93972700",
         463 => x"b387f900",
         464 => x"83a70700",
         465 => x"67800700",
         466 => x"9307f007",
         467 => x"630cf706",
         468 => x"6352640f",
         469 => x"9377f50f",
         470 => x"938607fe",
         471 => x"93f6f60f",
         472 => x"1306e005",
         473 => x"e36ed6fa",
         474 => x"b3868400",
         475 => x"2380f600",
         476 => x"13050700",
         477 => x"13041400",
         478 => x"ef008011",
         479 => x"6ff05ffa",
         480 => x"b3848400",
         481 => x"37150010",
         482 => x"23800400",
         483 => x"130505d9",
         484 => x"ef000012",
         485 => x"8320c102",
         486 => x"13050400",
         487 => x"03248102",
         488 => x"83244102",
         489 => x"03290102",
         490 => x"8329c101",
         491 => x"032a8101",
         492 => x"832a4101",
         493 => x"032b0101",
         494 => x"832bc100",
         495 => x"13010103",
         496 => x"67800000",
         497 => x"635a8002",
         498 => x"1305f007",
         499 => x"ef00400c",
         500 => x"1304f4ff",
         501 => x"6ff0dff4",
         502 => x"13854bd9",
         503 => x"ef00400d",
         504 => x"eff05fed",
         505 => x"1377f50f",
         506 => x"13040000",
         507 => x"e350e9f4",
         508 => x"9307f007",
         509 => x"e31ef7f4",
         510 => x"23248101",
         511 => x"130c5001",
         512 => x"13057000",
         513 => x"ef00c008",
         514 => x"eff0dfea",
         515 => x"1377f50f",
         516 => x"6348ec02",
         517 => x"032c8100",
         518 => x"6ff05ff1",
         519 => x"635a8002",
         520 => x"1305f007",
         521 => x"1304f4ff",
         522 => x"ef008006",
         523 => x"e31a04fe",
         524 => x"6ff01fef",
         525 => x"13057000",
         526 => x"ef008005",
         527 => x"6ff05fee",
         528 => x"9307f007",
         529 => x"e30ef7fa",
         530 => x"032c8100",
         531 => x"6ff05ff0",
         532 => x"eff05fe6",
         533 => x"1377f50f",
         534 => x"93075001",
         535 => x"e3d8e7ec",
         536 => x"6ff01ff9",
         537 => x"f32710fc",
         538 => x"63960700",
         539 => x"b7f7fa02",
         540 => x"93870708",
         541 => x"63060500",
         542 => x"33d5a702",
         543 => x"1305f5ff",
         544 => x"b70700f0",
         545 => x"23a6a702",
         546 => x"23a0b702",
         547 => x"67800000",
         548 => x"370700f0",
         549 => x"1375f50f",
         550 => x"13070702",
         551 => x"2324a700",
         552 => x"83274700",
         553 => x"93f70701",
         554 => x"e38c07fe",
         555 => x"67800000",
         556 => x"630e0502",
         557 => x"130101ff",
         558 => x"23248100",
         559 => x"23261100",
         560 => x"13040500",
         561 => x"03450500",
         562 => x"630a0500",
         563 => x"13041400",
         564 => x"eff01ffc",
         565 => x"03450400",
         566 => x"e31a05fe",
         567 => x"8320c100",
         568 => x"03248100",
         569 => x"13010101",
         570 => x"67800000",
         571 => x"67800000",
         572 => x"130101fe",
         573 => x"232e1100",
         574 => x"232c8100",
         575 => x"6350a00a",
         576 => x"23263101",
         577 => x"b7190010",
         578 => x"232a9100",
         579 => x"23282101",
         580 => x"23244101",
         581 => x"13090500",
         582 => x"93040000",
         583 => x"13040000",
         584 => x"9389d9c8",
         585 => x"130a1000",
         586 => x"6f000001",
         587 => x"3364c400",
         588 => x"93841400",
         589 => x"63029904",
         590 => x"eff0dfd7",
         591 => x"b387a900",
         592 => x"83c70700",
         593 => x"130605fd",
         594 => x"13144400",
         595 => x"13f74700",
         596 => x"93f64704",
         597 => x"e31c07fc",
         598 => x"93f73700",
         599 => x"e38a06fc",
         600 => x"63944701",
         601 => x"13050502",
         602 => x"130595fa",
         603 => x"93841400",
         604 => x"3364a400",
         605 => x"e31299fc",
         606 => x"8320c101",
         607 => x"13050400",
         608 => x"03248101",
         609 => x"83244101",
         610 => x"03290101",
         611 => x"8329c100",
         612 => x"032a8100",
         613 => x"13010102",
         614 => x"67800000",
         615 => x"13040000",
         616 => x"8320c101",
         617 => x"13050400",
         618 => x"03248101",
         619 => x"13010102",
         620 => x"67800000",
         621 => x"83470500",
         622 => x"37160010",
         623 => x"1306d6c8",
         624 => x"3307f600",
         625 => x"03470700",
         626 => x"93060500",
         627 => x"13758700",
         628 => x"630e0500",
         629 => x"83c71600",
         630 => x"93861600",
         631 => x"3307f600",
         632 => x"03470700",
         633 => x"13758700",
         634 => x"e31605fe",
         635 => x"13754704",
         636 => x"630a0506",
         637 => x"13050000",
         638 => x"13031000",
         639 => x"6f000002",
         640 => x"83c71600",
         641 => x"33e5a800",
         642 => x"93861600",
         643 => x"3307f600",
         644 => x"03470700",
         645 => x"13784704",
         646 => x"63000804",
         647 => x"13784700",
         648 => x"938807fd",
         649 => x"13773700",
         650 => x"13154500",
         651 => x"e31a08fc",
         652 => x"63146700",
         653 => x"93870702",
         654 => x"938797fa",
         655 => x"33e5a700",
         656 => x"83c71600",
         657 => x"93861600",
         658 => x"3307f600",
         659 => x"03470700",
         660 => x"13784704",
         661 => x"e31408fc",
         662 => x"63840500",
         663 => x"23a0d500",
         664 => x"67800000",
         665 => x"13050000",
         666 => x"6ff01fff",
         667 => x"130101fe",
         668 => x"232e1100",
         669 => x"23220100",
         670 => x"23240100",
         671 => x"23260100",
         672 => x"63040506",
         673 => x"232c8100",
         674 => x"93070500",
         675 => x"13040500",
         676 => x"63440504",
         677 => x"13074100",
         678 => x"1306a000",
         679 => x"13089000",
         680 => x"b3f6c702",
         681 => x"13050700",
         682 => x"1307f7ff",
         683 => x"93850700",
         684 => x"93860603",
         685 => x"a305d700",
         686 => x"b3d7c702",
         687 => x"e362b8fe",
         688 => x"3305c500",
         689 => x"eff0dfde",
         690 => x"8320c101",
         691 => x"03248101",
         692 => x"13010102",
         693 => x"67800000",
         694 => x"1305d002",
         695 => x"eff05fdb",
         696 => x"b3078040",
         697 => x"6ff01ffb",
         698 => x"13050003",
         699 => x"eff05fda",
         700 => x"8320c101",
         701 => x"13010102",
         702 => x"67800000",
         703 => x"130101fe",
         704 => x"232e1100",
         705 => x"23220100",
         706 => x"23240100",
         707 => x"23060100",
         708 => x"9387f5ff",
         709 => x"13077000",
         710 => x"6376f700",
         711 => x"93077000",
         712 => x"93058000",
         713 => x"13074100",
         714 => x"b307f700",
         715 => x"b385b740",
         716 => x"13069003",
         717 => x"9376f500",
         718 => x"13870603",
         719 => x"6374e600",
         720 => x"13877605",
         721 => x"2380e700",
         722 => x"9387f7ff",
         723 => x"13554500",
         724 => x"e392f5fe",
         725 => x"13054100",
         726 => x"eff09fd5",
         727 => x"8320c101",
         728 => x"13010102",
         729 => x"67800000",
         730 => x"130101ff",
         731 => x"23248100",
         732 => x"23229100",
         733 => x"37140010",
         734 => x"b7140010",
         735 => x"938784f1",
         736 => x"130484f1",
         737 => x"3304f440",
         738 => x"23202101",
         739 => x"23261100",
         740 => x"13542440",
         741 => x"938484f1",
         742 => x"13090000",
         743 => x"63108904",
         744 => x"b7140010",
         745 => x"37140010",
         746 => x"938784f1",
         747 => x"130484f1",
         748 => x"3304f440",
         749 => x"13542440",
         750 => x"938484f1",
         751 => x"13090000",
         752 => x"63188902",
         753 => x"8320c100",
         754 => x"03248100",
         755 => x"83244100",
         756 => x"03290100",
         757 => x"13010101",
         758 => x"67800000",
         759 => x"83a70400",
         760 => x"13091900",
         761 => x"93844400",
         762 => x"e7800700",
         763 => x"6ff01ffb",
         764 => x"83a70400",
         765 => x"13091900",
         766 => x"93844400",
         767 => x"e7800700",
         768 => x"6ff01ffc",
         769 => x"630a0602",
         770 => x"1306f6ff",
         771 => x"13070000",
         772 => x"b307e500",
         773 => x"b386e500",
         774 => x"83c70700",
         775 => x"83c60600",
         776 => x"6398d700",
         777 => x"6306c700",
         778 => x"13071700",
         779 => x"e39207fe",
         780 => x"3385d740",
         781 => x"67800000",
         782 => x"13050000",
         783 => x"67800000",
         784 => x"d8070010",
         785 => x"50070010",
         786 => x"50070010",
         787 => x"50070010",
         788 => x"50070010",
         789 => x"c4070010",
         790 => x"50070010",
         791 => x"80070010",
         792 => x"50070010",
         793 => x"50070010",
         794 => x"80070010",
         795 => x"50070010",
         796 => x"50070010",
         797 => x"50070010",
         798 => x"50070010",
         799 => x"50070010",
         800 => x"50070010",
         801 => x"50070010",
         802 => x"1c080010",
         803 => x"00202020",
         804 => x"20202020",
         805 => x"20202828",
         806 => x"28282820",
         807 => x"20202020",
         808 => x"20202020",
         809 => x"20202020",
         810 => x"20202020",
         811 => x"20881010",
         812 => x"10101010",
         813 => x"10101010",
         814 => x"10101010",
         815 => x"10040404",
         816 => x"04040404",
         817 => x"04040410",
         818 => x"10101010",
         819 => x"10104141",
         820 => x"41414141",
         821 => x"01010101",
         822 => x"01010101",
         823 => x"01010101",
         824 => x"01010101",
         825 => x"01010101",
         826 => x"10101010",
         827 => x"10104242",
         828 => x"42424242",
         829 => x"02020202",
         830 => x"02020202",
         831 => x"02020202",
         832 => x"02020202",
         833 => x"02020202",
         834 => x"10101010",
         835 => x"20000000",
         836 => x"00000000",
         837 => x"00000000",
         838 => x"00000000",
         839 => x"00000000",
         840 => x"00000000",
         841 => x"00000000",
         842 => x"00000000",
         843 => x"00000000",
         844 => x"00000000",
         845 => x"00000000",
         846 => x"00000000",
         847 => x"00000000",
         848 => x"00000000",
         849 => x"00000000",
         850 => x"00000000",
         851 => x"00000000",
         852 => x"00000000",
         853 => x"00000000",
         854 => x"00000000",
         855 => x"00000000",
         856 => x"00000000",
         857 => x"00000000",
         858 => x"00000000",
         859 => x"00000000",
         860 => x"00000000",
         861 => x"00000000",
         862 => x"00000000",
         863 => x"00000000",
         864 => x"00000000",
         865 => x"00000000",
         866 => x"00000000",
         867 => x"00000000",
         868 => x"0d0a0000",
         869 => x"3c627265",
         870 => x"616b3e0d",
         871 => x"0a000000",
         872 => x"54726170",
         873 => x"3a206d63",
         874 => x"61757365",
         875 => x"203d2030",
         876 => x"78000000",
         877 => x"0d0a5448",
         878 => x"55415320",
         879 => x"52495343",
         880 => x"2d562042",
         881 => x"6f6f746c",
         882 => x"6f616465",
         883 => x"72207630",
         884 => x"2e360d0a",
         885 => x"00000000",
         886 => x"436c6f63",
         887 => x"6b206672",
         888 => x"65717565",
         889 => x"6e63793a",
         890 => x"20000000",
         891 => x"3f0a0000",
         892 => x"3e200000",
         893 => x"68000000",
         894 => x"48656c70",
         895 => x"3a0d0a20",
         896 => x"68202020",
         897 => x"20202020",
         898 => x"20202020",
         899 => x"20202020",
         900 => x"202d2074",
         901 => x"68697320",
         902 => x"68656c70",
         903 => x"0d0a2072",
         904 => x"20202020",
         905 => x"20202020",
         906 => x"20202020",
         907 => x"20202020",
         908 => x"2d207275",
         909 => x"6e206170",
         910 => x"706c6963",
         911 => x"6174696f",
         912 => x"6e0d0a20",
         913 => x"7277203c",
         914 => x"61646472",
         915 => x"3e202020",
         916 => x"20202020",
         917 => x"202d2072",
         918 => x"65616420",
         919 => x"776f7264",
         920 => x"2066726f",
         921 => x"6d206164",
         922 => x"64720d0a",
         923 => x"20777720",
         924 => x"3c616464",
         925 => x"723e203c",
         926 => x"64617461",
         927 => x"3e202d20",
         928 => x"77726974",
         929 => x"6520776f",
         930 => x"72642064",
         931 => x"61746120",
         932 => x"61742061",
         933 => x"6464720d",
         934 => x"0a206477",
         935 => x"203c6164",
         936 => x"64723e20",
         937 => x"20202020",
         938 => x"2020202d",
         939 => x"2064756d",
         940 => x"70203136",
         941 => x"20776f72",
         942 => x"64730d0a",
         943 => x"206e2020",
         944 => x"20202020",
         945 => x"20202020",
         946 => x"20202020",
         947 => x"20202d20",
         948 => x"64756d70",
         949 => x"206e6578",
         950 => x"74203136",
         951 => x"20776f72",
         952 => x"64730000",
         953 => x"72000000",
         954 => x"72772000",
         955 => x"3a200000",
         956 => x"4e6f7420",
         957 => x"6f6e2034",
         958 => x"2d627974",
         959 => x"6520626f",
         960 => x"756e6461",
         961 => x"72792100",
         962 => x"77772000",
         963 => x"64772000",
         964 => x"20200000",
         965 => x"3f3f0000",
         966 => x"00000000"
            );
end package bootrom_image;
