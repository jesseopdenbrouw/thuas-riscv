-- #################################################################################################
-- # bootloader.vhd - The bootloader ROM                                                           #
-- # ********************************************************************************************* #
-- # This file is part of the THUAS RISCV RV32 Project                                             #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2023, Jesse op den Brouw. All rights reserved.                                  #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # https:/github.com/jesseopdenbrouw/riscv-rv32                                                  #
-- #################################################################################################

-- This file contains the description of the bootloader ROM. The ROM
-- is placed in immutable onboard RAM blocks. A read takes two
-- clock cycles, for both instruction and data.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.processor_common.all;

entity bootloader is
    generic (
          HAVE_BOOTLOADER_ROM : boolean
         );
    port (I_clk : in std_logic;
          I_areset : in std_logic;
          I_pc : in data_type;
          I_memaddress : in data_type;
          I_memsize : in memsize_type;
          I_csboot : in std_logic;
          I_stall : in std_logic;
          O_instr : out data_type;
          O_dataout : out data_type;
          O_memready : out std_logic;
          --
          O_load_misaligned_error : out std_logic
         );
end entity bootloader;

architecture rtl of bootloader is

-- The bootloader ROM
-- NOTE: the bootloader ROM is word (32 bits) size.
-- NOTE: data is in Little Endian format (as by the toolchain)
--       for half word and word entities
--       Set bootloader rom_size_bits as if it were bytes
--       default is 4 kB data
constant bootloader_size_bits : integer := 13;
constant bootloader_size : integer := 2**(bootloader_size_bits-2);
type bootloader_type is array(0 to bootloader_size-1) of data_type;

-- The bootloader ROM
signal bootrom : bootloader_type := (
           0 => x"97020000",
           1 => x"9382c207",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"9387c19a",
           8 => x"1387c185",
           9 => x"3386e740",
          10 => x"63f4e700",
          11 => x"13060000",
          12 => x"93050000",
          13 => x"1385c185",
          14 => x"ef008004",
          15 => x"37050020",
          16 => x"9387c185",
          17 => x"13070500",
          18 => x"3386e740",
          19 => x"63f4e700",
          20 => x"13060000",
          21 => x"b7250010",
          22 => x"938505e7",
          23 => x"13050500",
          24 => x"ef00c003",
          25 => x"ef10c048",
          26 => x"13060000",
          27 => x"9385c185",
          28 => x"13050000",
          29 => x"ef00c078",
          30 => x"ef00904b",
          31 => x"6f000000",
          32 => x"13030500",
          33 => x"630a0600",
          34 => x"2300b300",
          35 => x"1306f6ff",
          36 => x"13031300",
          37 => x"e31a06fe",
          38 => x"67800000",
          39 => x"13030500",
          40 => x"630e0600",
          41 => x"83830500",
          42 => x"23007300",
          43 => x"1306f6ff",
          44 => x"13031300",
          45 => x"93851500",
          46 => x"e31606fe",
          47 => x"67800000",
          48 => x"03460500",
          49 => x"83c60500",
          50 => x"13051500",
          51 => x"93851500",
          52 => x"6314d600",
          53 => x"e31606fe",
          54 => x"3305d640",
          55 => x"67800000",
          56 => x"6f000000",
          57 => x"13050000",
          58 => x"67800000",
          59 => x"13050000",
          60 => x"67800000",
          61 => x"130101ff",
          62 => x"23202101",
          63 => x"23261100",
          64 => x"13090600",
          65 => x"6356c002",
          66 => x"23248100",
          67 => x"23229100",
          68 => x"13840500",
          69 => x"b384c500",
          70 => x"03450400",
          71 => x"13041400",
          72 => x"eff05ffc",
          73 => x"e39a84fe",
          74 => x"03248100",
          75 => x"83244100",
          76 => x"8320c100",
          77 => x"13050900",
          78 => x"03290100",
          79 => x"13010101",
          80 => x"67800000",
          81 => x"130101ff",
          82 => x"23202101",
          83 => x"23261100",
          84 => x"13090600",
          85 => x"6356c002",
          86 => x"23248100",
          87 => x"23229100",
          88 => x"13840500",
          89 => x"b384c500",
          90 => x"eff05ff8",
          91 => x"13041400",
          92 => x"a30fa4fe",
          93 => x"e39a84fe",
          94 => x"03248100",
          95 => x"83244100",
          96 => x"8320c100",
          97 => x"13050900",
          98 => x"03290100",
          99 => x"13010101",
         100 => x"67800000",
         101 => x"13051000",
         102 => x"67800000",
         103 => x"130101ff",
         104 => x"23261100",
         105 => x"ef101020",
         106 => x"8320c100",
         107 => x"93076001",
         108 => x"2320f500",
         109 => x"1305f0ff",
         110 => x"13010101",
         111 => x"67800000",
         112 => x"1305f0ff",
         113 => x"67800000",
         114 => x"b7270000",
         115 => x"23a2f500",
         116 => x"13050000",
         117 => x"67800000",
         118 => x"13051000",
         119 => x"67800000",
         120 => x"13050000",
         121 => x"67800000",
         122 => x"130101fe",
         123 => x"2324c100",
         124 => x"2326d100",
         125 => x"2328e100",
         126 => x"232af100",
         127 => x"232c0101",
         128 => x"232e1101",
         129 => x"1305f0ff",
         130 => x"13010102",
         131 => x"67800000",
         132 => x"130101ff",
         133 => x"23261100",
         134 => x"ef10d018",
         135 => x"8320c100",
         136 => x"9307a000",
         137 => x"2320f500",
         138 => x"1305f0ff",
         139 => x"13010101",
         140 => x"67800000",
         141 => x"130101ff",
         142 => x"23261100",
         143 => x"ef109016",
         144 => x"8320c100",
         145 => x"93072000",
         146 => x"2320f500",
         147 => x"1305f0ff",
         148 => x"13010101",
         149 => x"67800000",
         150 => x"b7270000",
         151 => x"23a2f500",
         152 => x"13050000",
         153 => x"67800000",
         154 => x"130101ff",
         155 => x"23261100",
         156 => x"ef105013",
         157 => x"8320c100",
         158 => x"9307f001",
         159 => x"2320f500",
         160 => x"1305f0ff",
         161 => x"13010101",
         162 => x"67800000",
         163 => x"130101ff",
         164 => x"23261100",
         165 => x"ef101011",
         166 => x"8320c100",
         167 => x"9307b000",
         168 => x"2320f500",
         169 => x"1305f0ff",
         170 => x"13010101",
         171 => x"67800000",
         172 => x"130101ff",
         173 => x"23261100",
         174 => x"ef10d00e",
         175 => x"8320c100",
         176 => x"9307c000",
         177 => x"2320f500",
         178 => x"1305f0ff",
         179 => x"13010101",
         180 => x"67800000",
         181 => x"03a70186",
         182 => x"b7870020",
         183 => x"93870700",
         184 => x"93060040",
         185 => x"b387d740",
         186 => x"630c0700",
         187 => x"3305a700",
         188 => x"63e2a702",
         189 => x"23a0a186",
         190 => x"13050700",
         191 => x"67800000",
         192 => x"9386019b",
         193 => x"1387019b",
         194 => x"23a0d186",
         195 => x"3305a700",
         196 => x"e3f2a7fe",
         197 => x"130101ff",
         198 => x"23261100",
         199 => x"ef109008",
         200 => x"8320c100",
         201 => x"9307c000",
         202 => x"2320f500",
         203 => x"1307f0ff",
         204 => x"13050700",
         205 => x"13010101",
         206 => x"67800000",
         207 => x"b70700f0",
         208 => x"03a54702",
         209 => x"13754500",
         210 => x"67800000",
         211 => x"370700f0",
         212 => x"13070702",
         213 => x"83274700",
         214 => x"93f74700",
         215 => x"e38c07fe",
         216 => x"03258700",
         217 => x"1375f50f",
         218 => x"67800000",
         219 => x"130101fd",
         220 => x"232e3101",
         221 => x"b7290010",
         222 => x"23248102",
         223 => x"23229102",
         224 => x"23202103",
         225 => x"232c4101",
         226 => x"232a5101",
         227 => x"23286101",
         228 => x"23267101",
         229 => x"23261102",
         230 => x"93040500",
         231 => x"13040000",
         232 => x"9389c9ba",
         233 => x"13095001",
         234 => x"138bf5ff",
         235 => x"130a2000",
         236 => x"930a2001",
         237 => x"b72b0010",
         238 => x"eff05ff9",
         239 => x"1377f50f",
         240 => x"6340e902",
         241 => x"6352ea02",
         242 => x"9307d7ff",
         243 => x"63eefa00",
         244 => x"93972700",
         245 => x"b387f900",
         246 => x"83a70700",
         247 => x"67800700",
         248 => x"9307f007",
         249 => x"630cf706",
         250 => x"6352640f",
         251 => x"9377f50f",
         252 => x"938607fe",
         253 => x"93f6f60f",
         254 => x"1306e005",
         255 => x"e36ed6fa",
         256 => x"b3868400",
         257 => x"2380f600",
         258 => x"13050700",
         259 => x"13041400",
         260 => x"ef008011",
         261 => x"6ff05ffa",
         262 => x"b3848400",
         263 => x"37250010",
         264 => x"23800400",
         265 => x"130505c3",
         266 => x"ef000012",
         267 => x"8320c102",
         268 => x"13050400",
         269 => x"03248102",
         270 => x"83244102",
         271 => x"03290102",
         272 => x"8329c101",
         273 => x"032a8101",
         274 => x"832a4101",
         275 => x"032b0101",
         276 => x"832bc100",
         277 => x"13010103",
         278 => x"67800000",
         279 => x"635a8002",
         280 => x"1305f007",
         281 => x"ef00400c",
         282 => x"1304f4ff",
         283 => x"6ff0dff4",
         284 => x"13850bd6",
         285 => x"ef00400d",
         286 => x"eff05fed",
         287 => x"1377f50f",
         288 => x"13040000",
         289 => x"e350e9f4",
         290 => x"9307f007",
         291 => x"e31ef7f4",
         292 => x"23248101",
         293 => x"130c5001",
         294 => x"13057000",
         295 => x"ef00c008",
         296 => x"eff0dfea",
         297 => x"1377f50f",
         298 => x"6348ec02",
         299 => x"032c8100",
         300 => x"6ff05ff1",
         301 => x"635a8002",
         302 => x"1305f007",
         303 => x"1304f4ff",
         304 => x"ef008006",
         305 => x"e31a04fe",
         306 => x"6ff01fef",
         307 => x"13057000",
         308 => x"ef008005",
         309 => x"6ff05fee",
         310 => x"9307f007",
         311 => x"e30ef7fa",
         312 => x"032c8100",
         313 => x"6ff05ff0",
         314 => x"eff05fe6",
         315 => x"1377f50f",
         316 => x"93075001",
         317 => x"e3d8e7ec",
         318 => x"6ff01ff9",
         319 => x"f32710fc",
         320 => x"63960700",
         321 => x"b7f7fa02",
         322 => x"93870708",
         323 => x"63060500",
         324 => x"33d5a702",
         325 => x"1305f5ff",
         326 => x"b70700f0",
         327 => x"23a6a702",
         328 => x"23a0b702",
         329 => x"67800000",
         330 => x"370700f0",
         331 => x"1375f50f",
         332 => x"13070702",
         333 => x"2324a700",
         334 => x"83274700",
         335 => x"93f70701",
         336 => x"e38c07fe",
         337 => x"67800000",
         338 => x"630e0502",
         339 => x"130101ff",
         340 => x"23248100",
         341 => x"23261100",
         342 => x"13040500",
         343 => x"03450500",
         344 => x"630a0500",
         345 => x"13041400",
         346 => x"eff01ffc",
         347 => x"03450400",
         348 => x"e31a05fe",
         349 => x"8320c100",
         350 => x"03248100",
         351 => x"13010101",
         352 => x"67800000",
         353 => x"67800000",
         354 => x"130101fe",
         355 => x"232e1100",
         356 => x"232c8100",
         357 => x"6350a00a",
         358 => x"23263101",
         359 => x"b7290010",
         360 => x"232a9100",
         361 => x"23282101",
         362 => x"23244101",
         363 => x"13090500",
         364 => x"93040000",
         365 => x"13040000",
         366 => x"9389d9d6",
         367 => x"130a1000",
         368 => x"6f000001",
         369 => x"3364c400",
         370 => x"93841400",
         371 => x"63029904",
         372 => x"eff0dfd7",
         373 => x"b387a900",
         374 => x"83c70700",
         375 => x"130605fd",
         376 => x"13144400",
         377 => x"13f74700",
         378 => x"93f64704",
         379 => x"e31c07fc",
         380 => x"93f73700",
         381 => x"e38a06fc",
         382 => x"63944701",
         383 => x"13050502",
         384 => x"130595fa",
         385 => x"93841400",
         386 => x"3364a400",
         387 => x"e31299fc",
         388 => x"8320c101",
         389 => x"13050400",
         390 => x"03248101",
         391 => x"83244101",
         392 => x"03290101",
         393 => x"8329c100",
         394 => x"032a8100",
         395 => x"13010102",
         396 => x"67800000",
         397 => x"13040000",
         398 => x"8320c101",
         399 => x"13050400",
         400 => x"03248101",
         401 => x"13010102",
         402 => x"67800000",
         403 => x"83470500",
         404 => x"37260010",
         405 => x"1306d6d6",
         406 => x"3307f600",
         407 => x"03470700",
         408 => x"93060500",
         409 => x"13758700",
         410 => x"630e0500",
         411 => x"83c71600",
         412 => x"93861600",
         413 => x"3307f600",
         414 => x"03470700",
         415 => x"13758700",
         416 => x"e31605fe",
         417 => x"13754704",
         418 => x"630a0506",
         419 => x"13050000",
         420 => x"13031000",
         421 => x"6f000002",
         422 => x"83c71600",
         423 => x"33e5a800",
         424 => x"93861600",
         425 => x"3307f600",
         426 => x"03470700",
         427 => x"13784704",
         428 => x"63000804",
         429 => x"13784700",
         430 => x"938807fd",
         431 => x"13773700",
         432 => x"13154500",
         433 => x"e31a08fc",
         434 => x"63146700",
         435 => x"93870702",
         436 => x"938797fa",
         437 => x"33e5a700",
         438 => x"83c71600",
         439 => x"93861600",
         440 => x"3307f600",
         441 => x"03470700",
         442 => x"13784704",
         443 => x"e31408fc",
         444 => x"63840500",
         445 => x"23a0d500",
         446 => x"67800000",
         447 => x"13050000",
         448 => x"6ff01fff",
         449 => x"130101fe",
         450 => x"232e1100",
         451 => x"23220100",
         452 => x"23240100",
         453 => x"23260100",
         454 => x"63040506",
         455 => x"232c8100",
         456 => x"93070500",
         457 => x"13040500",
         458 => x"63440504",
         459 => x"13074100",
         460 => x"1306a000",
         461 => x"13089000",
         462 => x"b3f6c702",
         463 => x"13050700",
         464 => x"1307f7ff",
         465 => x"93850700",
         466 => x"93860603",
         467 => x"a305d700",
         468 => x"b3d7c702",
         469 => x"e362b8fe",
         470 => x"3305c500",
         471 => x"eff0dfde",
         472 => x"8320c101",
         473 => x"03248101",
         474 => x"13010102",
         475 => x"67800000",
         476 => x"1305d002",
         477 => x"eff05fdb",
         478 => x"b3078040",
         479 => x"6ff01ffb",
         480 => x"13050003",
         481 => x"eff05fda",
         482 => x"8320c101",
         483 => x"13010102",
         484 => x"67800000",
         485 => x"130101fe",
         486 => x"232e1100",
         487 => x"23220100",
         488 => x"23240100",
         489 => x"23060100",
         490 => x"9387f5ff",
         491 => x"13077000",
         492 => x"6376f700",
         493 => x"93077000",
         494 => x"93058000",
         495 => x"13074100",
         496 => x"b307f700",
         497 => x"b385b740",
         498 => x"13069003",
         499 => x"9376f500",
         500 => x"13870603",
         501 => x"6374e600",
         502 => x"13877605",
         503 => x"2380e700",
         504 => x"9387f7ff",
         505 => x"13554500",
         506 => x"e392f5fe",
         507 => x"13054100",
         508 => x"eff09fd5",
         509 => x"8320c101",
         510 => x"13010102",
         511 => x"67800000",
         512 => x"37c50100",
         513 => x"130101f8",
         514 => x"93050000",
         515 => x"13050520",
         516 => x"232e1106",
         517 => x"232c8106",
         518 => x"232a9106",
         519 => x"23282107",
         520 => x"23263107",
         521 => x"23244107",
         522 => x"23225107",
         523 => x"23206107",
         524 => x"232e7105",
         525 => x"232c8105",
         526 => x"232a9105",
         527 => x"2328a105",
         528 => x"2326b105",
         529 => x"eff09fcb",
         530 => x"37250010",
         531 => x"130585bf",
         532 => x"eff09fcf",
         533 => x"37250010",
         534 => x"1305c5c1",
         535 => x"eff0dfce",
         536 => x"732510fc",
         537 => x"37290010",
         538 => x"eff0dfe9",
         539 => x"130509c3",
         540 => x"eff09fcd",
         541 => x"b70700f0",
         542 => x"1307f03f",
         543 => x"370a1000",
         544 => x"b709a000",
         545 => x"23a2e700",
         546 => x"93041000",
         547 => x"130afaff",
         548 => x"b70a00f0",
         549 => x"93891900",
         550 => x"b3f74401",
         551 => x"639c0700",
         552 => x"1305a002",
         553 => x"eff05fc8",
         554 => x"83a74a00",
         555 => x"93d71700",
         556 => x"23a2fa00",
         557 => x"eff09fa8",
         558 => x"13040500",
         559 => x"63160504",
         560 => x"93841400",
         561 => x"e39a34fd",
         562 => x"b70700f0",
         563 => x"23a20700",
         564 => x"631a0400",
         565 => x"93050000",
         566 => x"13050000",
         567 => x"eff01fc2",
         568 => x"e7000400",
         569 => x"eff09fa6",
         570 => x"1375f50f",
         571 => x"93071002",
         572 => x"6300f502",
         573 => x"93074002",
         574 => x"93040000",
         575 => x"6316f520",
         576 => x"13041000",
         577 => x"6f00c001",
         578 => x"13041000",
         579 => x"6ff0dffb",
         580 => x"37250010",
         581 => x"130545c3",
         582 => x"eff01fc3",
         583 => x"13040000",
         584 => x"93040000",
         585 => x"370a00f0",
         586 => x"130b3005",
         587 => x"930ba004",
         588 => x"130c3002",
         589 => x"93092000",
         590 => x"930ca000",
         591 => x"b72a0010",
         592 => x"83274a00",
         593 => x"93c71700",
         594 => x"2322fa00",
         595 => x"eff01fa0",
         596 => x"1375f50f",
         597 => x"631e6517",
         598 => x"eff05f9f",
         599 => x"137df50f",
         600 => x"9307fdfc",
         601 => x"93f7f70f",
         602 => x"63e6f910",
         603 => x"93071003",
         604 => x"631afd04",
         605 => x"13052000",
         606 => x"eff01fc1",
         607 => x"930dd5ff",
         608 => x"13054000",
         609 => x"eff05fc0",
         610 => x"b70601ff",
         611 => x"b705ffff",
         612 => x"130d0500",
         613 => x"b38dad00",
         614 => x"9386f6ff",
         615 => x"9385f50f",
         616 => x"6318bd05",
         617 => x"130da000",
         618 => x"eff05f9a",
         619 => x"1375f50f",
         620 => x"e31ca5ff",
         621 => x"e31604f8",
         622 => x"13854ac3",
         623 => x"eff0dfb8",
         624 => x"6ff01ff8",
         625 => x"93072003",
         626 => x"13052000",
         627 => x"631afd00",
         628 => x"eff09fbb",
         629 => x"930dc5ff",
         630 => x"13056000",
         631 => x"6ff09ffa",
         632 => x"eff09fba",
         633 => x"930db5ff",
         634 => x"13058000",
         635 => x"6ff09ff9",
         636 => x"1378cdff",
         637 => x"13052000",
         638 => x"2326b100",
         639 => x"2324d100",
         640 => x"23220101",
         641 => x"eff05fb8",
         642 => x"03284100",
         643 => x"93070500",
         644 => x"37060001",
         645 => x"13753d00",
         646 => x"03270800",
         647 => x"83268100",
         648 => x"8325c100",
         649 => x"93083000",
         650 => x"1306f6ff",
         651 => x"13031000",
         652 => x"63063503",
         653 => x"630a1503",
         654 => x"630c6500",
         655 => x"137707f0",
         656 => x"b3e7e700",
         657 => x"2320f800",
         658 => x"130d1d00",
         659 => x"6ff05ff5",
         660 => x"3377b700",
         661 => x"93978700",
         662 => x"6ff09ffe",
         663 => x"3377d700",
         664 => x"93970701",
         665 => x"6ff0dffd",
         666 => x"3377c700",
         667 => x"93978701",
         668 => x"6ff01ffd",
         669 => x"93079dfc",
         670 => x"93f7f70f",
         671 => x"63e2f904",
         672 => x"13052000",
         673 => x"eff05fb0",
         674 => x"93077003",
         675 => x"13058000",
         676 => x"630afd00",
         677 => x"93078003",
         678 => x"13056000",
         679 => x"6304fd00",
         680 => x"13054000",
         681 => x"eff05fae",
         682 => x"93040500",
         683 => x"130da000",
         684 => x"eff0df89",
         685 => x"1375f50f",
         686 => x"e31ca5ff",
         687 => x"6ff09fef",
         688 => x"eff0df88",
         689 => x"1375f50f",
         690 => x"e31c95ff",
         691 => x"6ff09fee",
         692 => x"631e7509",
         693 => x"63180400",
         694 => x"37250010",
         695 => x"130545c3",
         696 => x"eff09fa6",
         697 => x"93050000",
         698 => x"13050000",
         699 => x"eff01fa1",
         700 => x"b70700f0",
         701 => x"23a20700",
         702 => x"e7800400",
         703 => x"b70700f0",
         704 => x"1307a00a",
         705 => x"23a2e700",
         706 => x"130509c3",
         707 => x"b7290010",
         708 => x"eff09fa3",
         709 => x"13040000",
         710 => x"372b0010",
         711 => x"b72b0010",
         712 => x"9389d9d6",
         713 => x"b7270010",
         714 => x"138587c3",
         715 => x"eff0dfa1",
         716 => x"93059002",
         717 => x"13054101",
         718 => x"eff05f83",
         719 => x"13054101",
         720 => x"ef00d024",
         721 => x"b7270010",
         722 => x"130a0500",
         723 => x"9385c7c3",
         724 => x"13054101",
         725 => x"eff0cfd6",
         726 => x"631e0500",
         727 => x"37250010",
         728 => x"130505c4",
         729 => x"eff05f9e",
         730 => x"6f004003",
         731 => x"e31485e5",
         732 => x"6ff0dff8",
         733 => x"b7270010",
         734 => x"9385c7d2",
         735 => x"13054101",
         736 => x"eff00fd4",
         737 => x"63100502",
         738 => x"93050000",
         739 => x"eff01f97",
         740 => x"b70700f0",
         741 => x"23a20700",
         742 => x"e7800400",
         743 => x"e3040af8",
         744 => x"6f004018",
         745 => x"b7270010",
         746 => x"13063000",
         747 => x"938507d3",
         748 => x"13054101",
         749 => x"ef000067",
         750 => x"63100504",
         751 => x"93050000",
         752 => x"13057101",
         753 => x"eff09fa8",
         754 => x"93773500",
         755 => x"13040500",
         756 => x"63940706",
         757 => x"93058000",
         758 => x"eff0dfbb",
         759 => x"37250010",
         760 => x"130545d3",
         761 => x"eff05f96",
         762 => x"03250400",
         763 => x"93058000",
         764 => x"eff05fba",
         765 => x"6ff09ffa",
         766 => x"13063000",
         767 => x"93050bd5",
         768 => x"13054101",
         769 => x"ef000062",
         770 => x"631e0502",
         771 => x"93050101",
         772 => x"13057101",
         773 => x"eff09fa3",
         774 => x"93773500",
         775 => x"13040500",
         776 => x"639c0700",
         777 => x"03250101",
         778 => x"93050000",
         779 => x"eff01fa2",
         780 => x"2320a400",
         781 => x"6ff09ff6",
         782 => x"37250010",
         783 => x"130585d3",
         784 => x"6ff05ff2",
         785 => x"13063000",
         786 => x"93854bd5",
         787 => x"13054101",
         788 => x"ef00405d",
         789 => x"83474101",
         790 => x"1307e006",
         791 => x"630c0508",
         792 => x"639ae70a",
         793 => x"93773400",
         794 => x"e39807fc",
         795 => x"130c0404",
         796 => x"b72c0010",
         797 => x"372d0010",
         798 => x"930d80ff",
         799 => x"93058000",
         800 => x"13050400",
         801 => x"eff01fb1",
         802 => x"13854cd3",
         803 => x"eff0df8b",
         804 => x"83270400",
         805 => x"93058000",
         806 => x"130a8001",
         807 => x"13850700",
         808 => x"2322f100",
         809 => x"eff01faf",
         810 => x"13058dd5",
         811 => x"eff0df89",
         812 => x"b70a00ff",
         813 => x"83274100",
         814 => x"33f55701",
         815 => x"33554501",
         816 => x"b3063501",
         817 => x"83c60600",
         818 => x"93f67609",
         819 => x"63800604",
         820 => x"130a8aff",
         821 => x"eff05f85",
         822 => x"93da8a00",
         823 => x"e31cbafd",
         824 => x"13044400",
         825 => x"130509c3",
         826 => x"eff01f86",
         827 => x"e31884f9",
         828 => x"6ff05fe3",
         829 => x"e388e7f6",
         830 => x"93050000",
         831 => x"13057101",
         832 => x"eff0df94",
         833 => x"13040500",
         834 => x"6ff0dff5",
         835 => x"1305e002",
         836 => x"6ff01ffc",
         837 => x"e3080ae0",
         838 => x"37250010",
         839 => x"1305c5d5",
         840 => x"eff09f82",
         841 => x"130509c3",
         842 => x"eff01f82",
         843 => x"6ff09fdf",
         844 => x"130101ff",
         845 => x"23248100",
         846 => x"23261100",
         847 => x"93070000",
         848 => x"13040500",
         849 => x"63880700",
         850 => x"93050000",
         851 => x"97000000",
         852 => x"e7000000",
         853 => x"83a74186",
         854 => x"63840700",
         855 => x"e7800700",
         856 => x"13050400",
         857 => x"eff0cfb7",
         858 => x"13050000",
         859 => x"67800000",
         860 => x"130101ff",
         861 => x"23248100",
         862 => x"23261100",
         863 => x"13040500",
         864 => x"2316b500",
         865 => x"2317c500",
         866 => x"23200500",
         867 => x"23220500",
         868 => x"23240500",
         869 => x"23220506",
         870 => x"23280500",
         871 => x"232a0500",
         872 => x"232c0500",
         873 => x"13068000",
         874 => x"93050000",
         875 => x"1305c505",
         876 => x"eff00fad",
         877 => x"b7170010",
         878 => x"9387870e",
         879 => x"2322f402",
         880 => x"b7170010",
         881 => x"93870714",
         882 => x"2324f402",
         883 => x"b7170010",
         884 => x"9387471c",
         885 => x"2326f402",
         886 => x"b7170010",
         887 => x"9387c721",
         888 => x"8320c100",
         889 => x"23208402",
         890 => x"2328f402",
         891 => x"03248100",
         892 => x"13010101",
         893 => x"67800000",
         894 => x"37060020",
         895 => x"b7250010",
         896 => x"37050020",
         897 => x"13060600",
         898 => x"938585ac",
         899 => x"1305c500",
         900 => x"6f008022",
         901 => x"83254500",
         902 => x"130101ff",
         903 => x"b7070020",
         904 => x"23248100",
         905 => x"23261100",
         906 => x"93874707",
         907 => x"13040500",
         908 => x"6384f500",
         909 => x"ef005049",
         910 => x"83258400",
         911 => x"9387c18d",
         912 => x"6386f500",
         913 => x"13050400",
         914 => x"ef001048",
         915 => x"8325c400",
         916 => x"93874194",
         917 => x"638cf500",
         918 => x"13050400",
         919 => x"03248100",
         920 => x"8320c100",
         921 => x"13010101",
         922 => x"6f001046",
         923 => x"8320c100",
         924 => x"03248100",
         925 => x"13010101",
         926 => x"67800000",
         927 => x"b7170010",
         928 => x"37050020",
         929 => x"130101ff",
         930 => x"938787df",
         931 => x"13060000",
         932 => x"93054000",
         933 => x"13054507",
         934 => x"23261100",
         935 => x"23a2f186",
         936 => x"eff01fed",
         937 => x"13061000",
         938 => x"93059000",
         939 => x"1385c18d",
         940 => x"eff01fec",
         941 => x"8320c100",
         942 => x"13062000",
         943 => x"93052001",
         944 => x"13854194",
         945 => x"13010101",
         946 => x"6ff09fea",
         947 => x"13050000",
         948 => x"67800000",
         949 => x"83a74186",
         950 => x"130101ff",
         951 => x"23202101",
         952 => x"23261100",
         953 => x"23248100",
         954 => x"23229100",
         955 => x"13090500",
         956 => x"63940700",
         957 => x"eff09ff8",
         958 => x"b7040020",
         959 => x"93840400",
         960 => x"03a48400",
         961 => x"83a74400",
         962 => x"9387f7ff",
         963 => x"63d80702",
         964 => x"83a70400",
         965 => x"6390070c",
         966 => x"9305c01a",
         967 => x"13050900",
         968 => x"ef005000",
         969 => x"13040500",
         970 => x"63140508",
         971 => x"23a00400",
         972 => x"9307c000",
         973 => x"2320f900",
         974 => x"6f004005",
         975 => x"0317c400",
         976 => x"63140706",
         977 => x"b707ffff",
         978 => x"93871700",
         979 => x"23220406",
         980 => x"23200400",
         981 => x"23220400",
         982 => x"23240400",
         983 => x"2326f400",
         984 => x"23280400",
         985 => x"232a0400",
         986 => x"232c0400",
         987 => x"13068000",
         988 => x"93050000",
         989 => x"1305c405",
         990 => x"eff08f90",
         991 => x"232a0402",
         992 => x"232c0402",
         993 => x"23240404",
         994 => x"23260404",
         995 => x"8320c100",
         996 => x"13050400",
         997 => x"03248100",
         998 => x"83244100",
         999 => x"03290100",
        1000 => x"13010101",
        1001 => x"67800000",
        1002 => x"13048406",
        1003 => x"6ff0dff5",
        1004 => x"93074000",
        1005 => x"23200500",
        1006 => x"2322f500",
        1007 => x"1305c500",
        1008 => x"2324a400",
        1009 => x"1306001a",
        1010 => x"93050000",
        1011 => x"eff04f8b",
        1012 => x"23a08400",
        1013 => x"83a40400",
        1014 => x"6ff09ff2",
        1015 => x"83270502",
        1016 => x"639e0700",
        1017 => x"b7170010",
        1018 => x"938747e1",
        1019 => x"2320f502",
        1020 => x"83a74186",
        1021 => x"63940700",
        1022 => x"6ff05fe8",
        1023 => x"67800000",
        1024 => x"67800000",
        1025 => x"67800000",
        1026 => x"37060020",
        1027 => x"b7150010",
        1028 => x"13060600",
        1029 => x"938585d6",
        1030 => x"13050000",
        1031 => x"6f00c001",
        1032 => x"37060020",
        1033 => x"b7150010",
        1034 => x"13060600",
        1035 => x"9385c5ec",
        1036 => x"13050000",
        1037 => x"6f004000",
        1038 => x"130101fd",
        1039 => x"23248102",
        1040 => x"23202103",
        1041 => x"232e3101",
        1042 => x"232c4101",
        1043 => x"23286101",
        1044 => x"23267101",
        1045 => x"23261102",
        1046 => x"23229102",
        1047 => x"232a5101",
        1048 => x"93090500",
        1049 => x"138a0500",
        1050 => x"13040600",
        1051 => x"13090000",
        1052 => x"130b1000",
        1053 => x"930bf0ff",
        1054 => x"83248400",
        1055 => x"832a4400",
        1056 => x"938afaff",
        1057 => x"63de0a02",
        1058 => x"03240400",
        1059 => x"e31604fe",
        1060 => x"8320c102",
        1061 => x"03248102",
        1062 => x"83244102",
        1063 => x"8329c101",
        1064 => x"032a8101",
        1065 => x"832a4101",
        1066 => x"032b0101",
        1067 => x"832bc100",
        1068 => x"13050900",
        1069 => x"03290102",
        1070 => x"13010103",
        1071 => x"67800000",
        1072 => x"83d7c400",
        1073 => x"637efb00",
        1074 => x"8397e400",
        1075 => x"638a7701",
        1076 => x"93850400",
        1077 => x"13850900",
        1078 => x"e7000a00",
        1079 => x"3369a900",
        1080 => x"93848406",
        1081 => x"6ff0dff9",
        1082 => x"130101ff",
        1083 => x"23248100",
        1084 => x"13840500",
        1085 => x"8395e500",
        1086 => x"23261100",
        1087 => x"ef004035",
        1088 => x"63400502",
        1089 => x"83274405",
        1090 => x"b387a700",
        1091 => x"232af404",
        1092 => x"8320c100",
        1093 => x"03248100",
        1094 => x"13010101",
        1095 => x"67800000",
        1096 => x"8357c400",
        1097 => x"37f7ffff",
        1098 => x"1307f7ff",
        1099 => x"b3f7e700",
        1100 => x"2316f400",
        1101 => x"6ff0dffd",
        1102 => x"13050000",
        1103 => x"67800000",
        1104 => x"83d7c500",
        1105 => x"130101fe",
        1106 => x"232c8100",
        1107 => x"232a9100",
        1108 => x"23282101",
        1109 => x"23263101",
        1110 => x"232e1100",
        1111 => x"93f70710",
        1112 => x"93040500",
        1113 => x"13840500",
        1114 => x"13090600",
        1115 => x"93890600",
        1116 => x"638a0700",
        1117 => x"8395e500",
        1118 => x"93062000",
        1119 => x"13060000",
        1120 => x"ef000028",
        1121 => x"8357c400",
        1122 => x"37f7ffff",
        1123 => x"1307f7ff",
        1124 => x"b3f7e700",
        1125 => x"8315e400",
        1126 => x"2316f400",
        1127 => x"03248101",
        1128 => x"8320c101",
        1129 => x"93860900",
        1130 => x"13060900",
        1131 => x"8329c100",
        1132 => x"03290101",
        1133 => x"13850400",
        1134 => x"83244101",
        1135 => x"13010102",
        1136 => x"6f00002e",
        1137 => x"130101ff",
        1138 => x"23248100",
        1139 => x"13840500",
        1140 => x"8395e500",
        1141 => x"23261100",
        1142 => x"ef008022",
        1143 => x"1307f0ff",
        1144 => x"8357c400",
        1145 => x"6312e502",
        1146 => x"37f7ffff",
        1147 => x"1307f7ff",
        1148 => x"b3f7e700",
        1149 => x"2316f400",
        1150 => x"8320c100",
        1151 => x"03248100",
        1152 => x"13010101",
        1153 => x"67800000",
        1154 => x"37170000",
        1155 => x"b3e7e700",
        1156 => x"2316f400",
        1157 => x"232aa404",
        1158 => x"6ff01ffe",
        1159 => x"8395e500",
        1160 => x"6f000004",
        1161 => x"630a0602",
        1162 => x"1306f6ff",
        1163 => x"13070000",
        1164 => x"b307e500",
        1165 => x"b386e500",
        1166 => x"83c70700",
        1167 => x"83c60600",
        1168 => x"6398d700",
        1169 => x"6306c700",
        1170 => x"13071700",
        1171 => x"e39207fe",
        1172 => x"3385d740",
        1173 => x"67800000",
        1174 => x"13050000",
        1175 => x"67800000",
        1176 => x"130101ff",
        1177 => x"23248100",
        1178 => x"23229100",
        1179 => x"13040500",
        1180 => x"13850500",
        1181 => x"23261100",
        1182 => x"23a40186",
        1183 => x"efe05ff4",
        1184 => x"9307f0ff",
        1185 => x"6318f500",
        1186 => x"83a78186",
        1187 => x"63840700",
        1188 => x"2320f400",
        1189 => x"8320c100",
        1190 => x"03248100",
        1191 => x"83244100",
        1192 => x"13010101",
        1193 => x"67800000",
        1194 => x"83a78185",
        1195 => x"6388a714",
        1196 => x"8327c501",
        1197 => x"130101fe",
        1198 => x"232c8100",
        1199 => x"232e1100",
        1200 => x"232a9100",
        1201 => x"23282101",
        1202 => x"23263101",
        1203 => x"13040500",
        1204 => x"638a0704",
        1205 => x"83a7c700",
        1206 => x"638c0702",
        1207 => x"93040000",
        1208 => x"13090008",
        1209 => x"8327c401",
        1210 => x"83a7c700",
        1211 => x"b3879700",
        1212 => x"83a50700",
        1213 => x"639c050c",
        1214 => x"93844400",
        1215 => x"e39424ff",
        1216 => x"8327c401",
        1217 => x"13050400",
        1218 => x"83a5c700",
        1219 => x"ef00c029",
        1220 => x"8327c401",
        1221 => x"83a50700",
        1222 => x"63860500",
        1223 => x"13050400",
        1224 => x"ef008028",
        1225 => x"83254401",
        1226 => x"63860500",
        1227 => x"13050400",
        1228 => x"ef008027",
        1229 => x"8325c401",
        1230 => x"63860500",
        1231 => x"13050400",
        1232 => x"ef008026",
        1233 => x"83250403",
        1234 => x"63860500",
        1235 => x"13050400",
        1236 => x"ef008025",
        1237 => x"83254403",
        1238 => x"63860500",
        1239 => x"13050400",
        1240 => x"ef008024",
        1241 => x"83258403",
        1242 => x"63860500",
        1243 => x"13050400",
        1244 => x"ef008023",
        1245 => x"83258404",
        1246 => x"63860500",
        1247 => x"13050400",
        1248 => x"ef008022",
        1249 => x"83254404",
        1250 => x"63860500",
        1251 => x"13050400",
        1252 => x"ef008021",
        1253 => x"8325c402",
        1254 => x"63860500",
        1255 => x"13050400",
        1256 => x"ef008020",
        1257 => x"83270402",
        1258 => x"638c0702",
        1259 => x"13050400",
        1260 => x"03248101",
        1261 => x"8320c101",
        1262 => x"83244101",
        1263 => x"03290101",
        1264 => x"8329c100",
        1265 => x"13010102",
        1266 => x"67800700",
        1267 => x"83a90500",
        1268 => x"13050400",
        1269 => x"ef00401d",
        1270 => x"93850900",
        1271 => x"6ff09ff1",
        1272 => x"8320c101",
        1273 => x"03248101",
        1274 => x"83244101",
        1275 => x"03290101",
        1276 => x"8329c100",
        1277 => x"13010102",
        1278 => x"67800000",
        1279 => x"67800000",
        1280 => x"130101ff",
        1281 => x"23248100",
        1282 => x"23229100",
        1283 => x"13040500",
        1284 => x"13850500",
        1285 => x"93050600",
        1286 => x"13860600",
        1287 => x"23261100",
        1288 => x"23a40186",
        1289 => x"efe0dfdb",
        1290 => x"9307f0ff",
        1291 => x"6318f500",
        1292 => x"83a78186",
        1293 => x"63840700",
        1294 => x"2320f400",
        1295 => x"8320c100",
        1296 => x"03248100",
        1297 => x"83244100",
        1298 => x"13010101",
        1299 => x"67800000",
        1300 => x"130101ff",
        1301 => x"23248100",
        1302 => x"23229100",
        1303 => x"13040500",
        1304 => x"13850500",
        1305 => x"93050600",
        1306 => x"13860600",
        1307 => x"23261100",
        1308 => x"23a40186",
        1309 => x"efe01fcd",
        1310 => x"9307f0ff",
        1311 => x"6318f500",
        1312 => x"83a78186",
        1313 => x"63840700",
        1314 => x"2320f400",
        1315 => x"8320c100",
        1316 => x"03248100",
        1317 => x"83244100",
        1318 => x"13010101",
        1319 => x"67800000",
        1320 => x"130101ff",
        1321 => x"23248100",
        1322 => x"23229100",
        1323 => x"13040500",
        1324 => x"13850500",
        1325 => x"93050600",
        1326 => x"13860600",
        1327 => x"23261100",
        1328 => x"23a40186",
        1329 => x"efe01fc3",
        1330 => x"9307f0ff",
        1331 => x"6318f500",
        1332 => x"83a78186",
        1333 => x"63840700",
        1334 => x"2320f400",
        1335 => x"8320c100",
        1336 => x"03248100",
        1337 => x"83244100",
        1338 => x"13010101",
        1339 => x"67800000",
        1340 => x"130101ff",
        1341 => x"23248100",
        1342 => x"23229100",
        1343 => x"37240010",
        1344 => x"b7240010",
        1345 => x"938704e7",
        1346 => x"130404e7",
        1347 => x"3304f440",
        1348 => x"23202101",
        1349 => x"23261100",
        1350 => x"13542440",
        1351 => x"938404e7",
        1352 => x"13090000",
        1353 => x"63108904",
        1354 => x"b7240010",
        1355 => x"37240010",
        1356 => x"938704e7",
        1357 => x"130404e7",
        1358 => x"3304f440",
        1359 => x"13542440",
        1360 => x"938404e7",
        1361 => x"13090000",
        1362 => x"63188902",
        1363 => x"8320c100",
        1364 => x"03248100",
        1365 => x"83244100",
        1366 => x"03290100",
        1367 => x"13010101",
        1368 => x"67800000",
        1369 => x"83a70400",
        1370 => x"13091900",
        1371 => x"93844400",
        1372 => x"e7800700",
        1373 => x"6ff01ffb",
        1374 => x"83a70400",
        1375 => x"13091900",
        1376 => x"93844400",
        1377 => x"e7800700",
        1378 => x"6ff01ffc",
        1379 => x"93070500",
        1380 => x"03c70700",
        1381 => x"93871700",
        1382 => x"e31c07fe",
        1383 => x"3385a740",
        1384 => x"1305f5ff",
        1385 => x"67800000",
        1386 => x"638a050e",
        1387 => x"83a7c5ff",
        1388 => x"130101fe",
        1389 => x"232c8100",
        1390 => x"232e1100",
        1391 => x"1384c5ff",
        1392 => x"63d40700",
        1393 => x"3304f400",
        1394 => x"2326a100",
        1395 => x"ef008031",
        1396 => x"83a70187",
        1397 => x"0325c100",
        1398 => x"639e0700",
        1399 => x"23220400",
        1400 => x"23a88186",
        1401 => x"03248101",
        1402 => x"8320c101",
        1403 => x"13010102",
        1404 => x"6f00802f",
        1405 => x"6374f402",
        1406 => x"03260400",
        1407 => x"b306c400",
        1408 => x"639ad700",
        1409 => x"83a60700",
        1410 => x"83a74700",
        1411 => x"b386c600",
        1412 => x"2320d400",
        1413 => x"2322f400",
        1414 => x"6ff09ffc",
        1415 => x"13870700",
        1416 => x"83a74700",
        1417 => x"63840700",
        1418 => x"e37af4fe",
        1419 => x"83260700",
        1420 => x"3306d700",
        1421 => x"63188602",
        1422 => x"03260400",
        1423 => x"b386c600",
        1424 => x"2320d700",
        1425 => x"3306d700",
        1426 => x"e39ec7f8",
        1427 => x"03a60700",
        1428 => x"83a74700",
        1429 => x"b306d600",
        1430 => x"2320d700",
        1431 => x"2322f700",
        1432 => x"6ff05ff8",
        1433 => x"6378c400",
        1434 => x"9307c000",
        1435 => x"2320f500",
        1436 => x"6ff05ff7",
        1437 => x"03260400",
        1438 => x"b306c400",
        1439 => x"639ad700",
        1440 => x"83a60700",
        1441 => x"83a74700",
        1442 => x"b386c600",
        1443 => x"2320d400",
        1444 => x"2322f400",
        1445 => x"23228700",
        1446 => x"6ff0dff4",
        1447 => x"67800000",
        1448 => x"130101ff",
        1449 => x"23202101",
        1450 => x"83a7c186",
        1451 => x"23248100",
        1452 => x"23229100",
        1453 => x"23261100",
        1454 => x"93040500",
        1455 => x"13840500",
        1456 => x"63980700",
        1457 => x"93050000",
        1458 => x"ef004049",
        1459 => x"23a6a186",
        1460 => x"93050400",
        1461 => x"13850400",
        1462 => x"ef004048",
        1463 => x"1309f0ff",
        1464 => x"63122503",
        1465 => x"1304f0ff",
        1466 => x"8320c100",
        1467 => x"13050400",
        1468 => x"03248100",
        1469 => x"83244100",
        1470 => x"03290100",
        1471 => x"13010101",
        1472 => x"67800000",
        1473 => x"13043500",
        1474 => x"1374c4ff",
        1475 => x"e30e85fc",
        1476 => x"b305a440",
        1477 => x"13850400",
        1478 => x"ef004044",
        1479 => x"e31625fd",
        1480 => x"6ff05ffc",
        1481 => x"130101fe",
        1482 => x"232a9100",
        1483 => x"93843500",
        1484 => x"93f4c4ff",
        1485 => x"23282101",
        1486 => x"232e1100",
        1487 => x"232c8100",
        1488 => x"23263101",
        1489 => x"23244101",
        1490 => x"93848400",
        1491 => x"9307c000",
        1492 => x"13090500",
        1493 => x"63f0f40a",
        1494 => x"9304c000",
        1495 => x"63eeb408",
        1496 => x"13050900",
        1497 => x"ef000018",
        1498 => x"83a70187",
        1499 => x"13840700",
        1500 => x"631a040a",
        1501 => x"93850400",
        1502 => x"13050900",
        1503 => x"eff05ff2",
        1504 => x"9307f0ff",
        1505 => x"13040500",
        1506 => x"6316f514",
        1507 => x"03a40187",
        1508 => x"93070400",
        1509 => x"639c0710",
        1510 => x"63040412",
        1511 => x"032a0400",
        1512 => x"93050000",
        1513 => x"13050900",
        1514 => x"330a4401",
        1515 => x"ef00003b",
        1516 => x"6318aa10",
        1517 => x"83270400",
        1518 => x"13050900",
        1519 => x"b384f440",
        1520 => x"93850400",
        1521 => x"eff0dfed",
        1522 => x"9307f0ff",
        1523 => x"630af50e",
        1524 => x"83270400",
        1525 => x"b3879700",
        1526 => x"2320f400",
        1527 => x"83a70187",
        1528 => x"638e070e",
        1529 => x"03a74700",
        1530 => x"6318870c",
        1531 => x"23a20700",
        1532 => x"6f004006",
        1533 => x"e3d404f6",
        1534 => x"9307c000",
        1535 => x"2320f900",
        1536 => x"13050000",
        1537 => x"8320c101",
        1538 => x"03248101",
        1539 => x"83244101",
        1540 => x"03290101",
        1541 => x"8329c100",
        1542 => x"032a8100",
        1543 => x"13010102",
        1544 => x"67800000",
        1545 => x"83260400",
        1546 => x"b3869640",
        1547 => x"63ca0606",
        1548 => x"1307b000",
        1549 => x"637ad704",
        1550 => x"23209400",
        1551 => x"33079400",
        1552 => x"63908704",
        1553 => x"23a8e186",
        1554 => x"83274400",
        1555 => x"2320d700",
        1556 => x"2322f700",
        1557 => x"13050900",
        1558 => x"ef000009",
        1559 => x"1305b400",
        1560 => x"93074400",
        1561 => x"137585ff",
        1562 => x"3307f540",
        1563 => x"e30cf5f8",
        1564 => x"3304e400",
        1565 => x"b387a740",
        1566 => x"2320f400",
        1567 => x"6ff09ff8",
        1568 => x"23a2e700",
        1569 => x"6ff05ffc",
        1570 => x"03274400",
        1571 => x"63968700",
        1572 => x"23a8e186",
        1573 => x"6ff01ffc",
        1574 => x"23a2e700",
        1575 => x"6ff09ffb",
        1576 => x"93070400",
        1577 => x"03244400",
        1578 => x"6ff09fec",
        1579 => x"13840700",
        1580 => x"83a74700",
        1581 => x"6ff01fee",
        1582 => x"93070700",
        1583 => x"6ff05ff2",
        1584 => x"9307c000",
        1585 => x"2320f900",
        1586 => x"13050900",
        1587 => x"ef00c001",
        1588 => x"6ff01ff3",
        1589 => x"23209500",
        1590 => x"6ff0dff7",
        1591 => x"23220000",
        1592 => x"73001000",
        1593 => x"67800000",
        1594 => x"67800000",
        1595 => x"8397c500",
        1596 => x"130101fe",
        1597 => x"232c8100",
        1598 => x"232a9100",
        1599 => x"232e1100",
        1600 => x"23282101",
        1601 => x"23263101",
        1602 => x"13f78700",
        1603 => x"93040500",
        1604 => x"13840500",
        1605 => x"631a0712",
        1606 => x"03a74500",
        1607 => x"6346e000",
        1608 => x"03a70504",
        1609 => x"6356e010",
        1610 => x"0327c402",
        1611 => x"63020710",
        1612 => x"03a90400",
        1613 => x"93963701",
        1614 => x"23a00400",
        1615 => x"83250402",
        1616 => x"63dc060a",
        1617 => x"03264405",
        1618 => x"8357c400",
        1619 => x"93f74700",
        1620 => x"638e0700",
        1621 => x"83274400",
        1622 => x"3306f640",
        1623 => x"83274403",
        1624 => x"63860700",
        1625 => x"83270404",
        1626 => x"3306f640",
        1627 => x"8327c402",
        1628 => x"83250402",
        1629 => x"93060000",
        1630 => x"13850400",
        1631 => x"e7800700",
        1632 => x"1307f0ff",
        1633 => x"8357c400",
        1634 => x"6312e502",
        1635 => x"83a60400",
        1636 => x"1307d001",
        1637 => x"6362d70a",
        1638 => x"37074020",
        1639 => x"13071700",
        1640 => x"3357d700",
        1641 => x"13771700",
        1642 => x"63080708",
        1643 => x"03270401",
        1644 => x"23220400",
        1645 => x"2320e400",
        1646 => x"13973701",
        1647 => x"635c0700",
        1648 => x"9307f0ff",
        1649 => x"6316f500",
        1650 => x"83a70400",
        1651 => x"63940700",
        1652 => x"232aa404",
        1653 => x"83254403",
        1654 => x"23a02401",
        1655 => x"638a0504",
        1656 => x"93074404",
        1657 => x"6386f500",
        1658 => x"13850400",
        1659 => x"eff0dfbb",
        1660 => x"232a0402",
        1661 => x"6f00c003",
        1662 => x"13060000",
        1663 => x"93061000",
        1664 => x"13850400",
        1665 => x"e7000700",
        1666 => x"9307f0ff",
        1667 => x"13060500",
        1668 => x"e31cf5f2",
        1669 => x"83a70400",
        1670 => x"e38807f2",
        1671 => x"1307d001",
        1672 => x"6386e700",
        1673 => x"13076001",
        1674 => x"6394e706",
        1675 => x"23a02401",
        1676 => x"13050000",
        1677 => x"6f00c006",
        1678 => x"93e70704",
        1679 => x"93970701",
        1680 => x"93d70741",
        1681 => x"6f004005",
        1682 => x"83a90501",
        1683 => x"e38209fe",
        1684 => x"03a90500",
        1685 => x"93f73700",
        1686 => x"23a03501",
        1687 => x"33093941",
        1688 => x"13070000",
        1689 => x"63940700",
        1690 => x"03a74501",
        1691 => x"2324e400",
        1692 => x"e35020fd",
        1693 => x"83278402",
        1694 => x"83250402",
        1695 => x"93060900",
        1696 => x"13860900",
        1697 => x"13850400",
        1698 => x"e7800700",
        1699 => x"6348a002",
        1700 => x"8317c400",
        1701 => x"93e70704",
        1702 => x"2316f400",
        1703 => x"1305f0ff",
        1704 => x"8320c101",
        1705 => x"03248101",
        1706 => x"83244101",
        1707 => x"03290101",
        1708 => x"8329c100",
        1709 => x"13010102",
        1710 => x"67800000",
        1711 => x"b389a900",
        1712 => x"3309a940",
        1713 => x"6ff0dffa",
        1714 => x"83a70501",
        1715 => x"638e0704",
        1716 => x"130101fe",
        1717 => x"232c8100",
        1718 => x"232e1100",
        1719 => x"13040500",
        1720 => x"630c0500",
        1721 => x"83270502",
        1722 => x"63980700",
        1723 => x"2326b100",
        1724 => x"eff0cfce",
        1725 => x"8325c100",
        1726 => x"8397c500",
        1727 => x"638c0700",
        1728 => x"13050400",
        1729 => x"03248101",
        1730 => x"8320c101",
        1731 => x"13010102",
        1732 => x"6ff0dfdd",
        1733 => x"8320c101",
        1734 => x"03248101",
        1735 => x"13050000",
        1736 => x"13010102",
        1737 => x"67800000",
        1738 => x"13050000",
        1739 => x"67800000",
        1740 => x"93050500",
        1741 => x"63100502",
        1742 => x"37060020",
        1743 => x"b7250010",
        1744 => x"37050020",
        1745 => x"13060600",
        1746 => x"938585ac",
        1747 => x"1305c500",
        1748 => x"6ff08fce",
        1749 => x"03a58185",
        1750 => x"6ff01ff7",
        1751 => x"130101ff",
        1752 => x"23248100",
        1753 => x"23229100",
        1754 => x"13040500",
        1755 => x"13850500",
        1756 => x"23261100",
        1757 => x"23a40186",
        1758 => x"efe0cff5",
        1759 => x"9307f0ff",
        1760 => x"6318f500",
        1761 => x"83a78186",
        1762 => x"63840700",
        1763 => x"2320f400",
        1764 => x"8320c100",
        1765 => x"03248100",
        1766 => x"83244100",
        1767 => x"13010101",
        1768 => x"67800000",
        1769 => x"03a58185",
        1770 => x"67800000",
        1771 => x"70040010",
        1772 => x"e8030010",
        1773 => x"e8030010",
        1774 => x"e8030010",
        1775 => x"e8030010",
        1776 => x"5c040010",
        1777 => x"e8030010",
        1778 => x"18040010",
        1779 => x"e8030010",
        1780 => x"e8030010",
        1781 => x"18040010",
        1782 => x"e8030010",
        1783 => x"e8030010",
        1784 => x"e8030010",
        1785 => x"e8030010",
        1786 => x"e8030010",
        1787 => x"e8030010",
        1788 => x"e8030010",
        1789 => x"b4040010",
        1790 => x"0d0a5448",
        1791 => x"55415320",
        1792 => x"52495343",
        1793 => x"2d562042",
        1794 => x"6f6f746c",
        1795 => x"6f616465",
        1796 => x"72207630",
        1797 => x"2e350d0a",
        1798 => x"00000000",
        1799 => x"436c6f63",
        1800 => x"6b206672",
        1801 => x"65717565",
        1802 => x"6e63793a",
        1803 => x"20000000",
        1804 => x"0d0a0000",
        1805 => x"3f0a0000",
        1806 => x"3e200000",
        1807 => x"68000000",
        1808 => x"48656c70",
        1809 => x"3a0d0a20",
        1810 => x"68202020",
        1811 => x"20202020",
        1812 => x"20202020",
        1813 => x"20202020",
        1814 => x"202d2074",
        1815 => x"68697320",
        1816 => x"68656c70",
        1817 => x"0d0a2072",
        1818 => x"20202020",
        1819 => x"20202020",
        1820 => x"20202020",
        1821 => x"20202020",
        1822 => x"2d207275",
        1823 => x"6e206170",
        1824 => x"706c6963",
        1825 => x"6174696f",
        1826 => x"6e0d0a20",
        1827 => x"7277203c",
        1828 => x"61646472",
        1829 => x"3e202020",
        1830 => x"20202020",
        1831 => x"202d2072",
        1832 => x"65616420",
        1833 => x"776f7264",
        1834 => x"2066726f",
        1835 => x"6d206164",
        1836 => x"64720d0a",
        1837 => x"20777720",
        1838 => x"3c616464",
        1839 => x"723e203c",
        1840 => x"64617461",
        1841 => x"3e202d20",
        1842 => x"77726974",
        1843 => x"6520776f",
        1844 => x"72642064",
        1845 => x"61746120",
        1846 => x"61742061",
        1847 => x"6464720d",
        1848 => x"0a206477",
        1849 => x"203c6164",
        1850 => x"64723e20",
        1851 => x"20202020",
        1852 => x"2020202d",
        1853 => x"2064756d",
        1854 => x"70203136",
        1855 => x"20776f72",
        1856 => x"64730d0a",
        1857 => x"206e2020",
        1858 => x"20202020",
        1859 => x"20202020",
        1860 => x"20202020",
        1861 => x"20202d20",
        1862 => x"64756d70",
        1863 => x"206e6578",
        1864 => x"74203136",
        1865 => x"20776f72",
        1866 => x"64730000",
        1867 => x"72000000",
        1868 => x"72772000",
        1869 => x"3a200000",
        1870 => x"4e6f7420",
        1871 => x"6f6e2034",
        1872 => x"2d627974",
        1873 => x"6520626f",
        1874 => x"756e6461",
        1875 => x"72792100",
        1876 => x"77772000",
        1877 => x"64772000",
        1878 => x"20200000",
        1879 => x"3f3f0000",
        1880 => x"3c627265",
        1881 => x"616b3e0d",
        1882 => x"0a000000",
        1883 => x"00202020",
        1884 => x"20202020",
        1885 => x"20202828",
        1886 => x"28282820",
        1887 => x"20202020",
        1888 => x"20202020",
        1889 => x"20202020",
        1890 => x"20202020",
        1891 => x"20881010",
        1892 => x"10101010",
        1893 => x"10101010",
        1894 => x"10101010",
        1895 => x"10040404",
        1896 => x"04040404",
        1897 => x"04040410",
        1898 => x"10101010",
        1899 => x"10104141",
        1900 => x"41414141",
        1901 => x"01010101",
        1902 => x"01010101",
        1903 => x"01010101",
        1904 => x"01010101",
        1905 => x"01010101",
        1906 => x"10101010",
        1907 => x"10104242",
        1908 => x"42424242",
        1909 => x"02020202",
        1910 => x"02020202",
        1911 => x"02020202",
        1912 => x"02020202",
        1913 => x"02020202",
        1914 => x"10101010",
        1915 => x"20000000",
        1916 => x"00000000",
        1917 => x"00000000",
        1918 => x"00000000",
        1919 => x"00000000",
        1920 => x"00000000",
        1921 => x"00000000",
        1922 => x"00000000",
        1923 => x"00000000",
        1924 => x"00000000",
        1925 => x"00000000",
        1926 => x"00000000",
        1927 => x"00000000",
        1928 => x"00000000",
        1929 => x"00000000",
        1930 => x"00000000",
        1931 => x"00000000",
        1932 => x"00000000",
        1933 => x"00000000",
        1934 => x"00000000",
        1935 => x"00000000",
        1936 => x"00000000",
        1937 => x"00000000",
        1938 => x"00000000",
        1939 => x"00000000",
        1940 => x"00000000",
        1941 => x"00000000",
        1942 => x"00000000",
        1943 => x"00000000",
        1944 => x"00000000",
        1945 => x"00000000",
        1946 => x"00000000",
        1947 => x"00000000",
        1948 => x"00000000",
        1949 => x"03000000",
        1950 => x"74000020",
        1951 => x"00000000",
        1952 => x"74000020",
        1953 => x"dc000020",
        1954 => x"44010020",
        1955 => x"00000000",
        1956 => x"00000000",
        1957 => x"00000000",
        1958 => x"00000000",
        1959 => x"00000000",
        1960 => x"00000000",
        1961 => x"00000000",
        1962 => x"00000000",
        1963 => x"00000000",
        1964 => x"00000000",
        1965 => x"00000000",
        1966 => x"00000000",
        1967 => x"00000000",
        1968 => x"00000000",
        1969 => x"00000000",
        1970 => x"0c000020",
         others => (others => '0')
        );

begin

    gen_bootrom: if HAVE_BOOTLOADER_ROM generate

        -- Boot ROM, for both instructions and read-only data
        process (I_clk, I_areset, I_pc, I_memaddress, I_csboot, I_memsize, I_stall) is
        variable address_instr : integer range 0 to bootloader_size-1;
        variable address_data : integer range 0 to bootloader_size-1;
        variable instr_var : data_type;
        variable instr_recode : data_type;
        variable romdata_var : data_type;
        constant x : data_type := (others => 'X');
        begin
            -- Calculate addresses
            address_instr := to_integer(unsigned(I_pc(bootloader_size_bits-1 downto 2)));
            address_data := to_integer(unsigned(I_memaddress(bootloader_size_bits-1 downto 2)));

            -- Quartus will detect ROM table and uses onboard RAM
            -- Do not use reset, otherwise ROM will be created with ALMs
            if rising_edge(I_clk) then
                if I_stall = '0' then
                    instr_var := bootrom(address_instr);
                end if;
                romdata_var := bootrom(address_data);
            end if;
            
            -- Recode instruction
            O_instr <= instr_var(7 downto 0) & instr_var(15 downto 8) & instr_var(23 downto 16) & instr_var(31 downto 24);
            
            O_load_misaligned_error <= '0';
            
            -- By natural size, for data
            if I_csboot = '1' then
                if I_memsize = memsize_word and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= romdata_var(7 downto 0) & romdata_var(15 downto 8) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= x(31 downto 16) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "10" then
                    O_dataout <= x(31 downto 16) & romdata_var(7 downto 0) & romdata_var(15 downto 8);
                elsif I_memsize = memsize_byte then
                    case I_memaddress(1 downto 0) is
                        when "00" => O_dataout <= x(31 downto 8) & romdata_var(31 downto 24);
                        when "01" => O_dataout <= x(31 downto 8) & romdata_var(23 downto 16);
                        when "10" => O_dataout <= x(31 downto 8) & romdata_var(15 downto 8);
                        when "11" => O_dataout <= x(31 downto 8) & romdata_var(7 downto 0);
                        when others => O_dataout <= x; O_load_misaligned_error <= '1';
                    end case;
                else
                    -- Chip select, but not aligned
                    O_dataout <= x;
                    O_load_misaligned_error <= '1';
                end if;
            else
                -- No chip select, so no data
                O_dataout <= x;
            end if;
        end process;
        
        -- Generate boot ROM ready signal for reads and writes    
        process (I_clk, I_areset, I_csboot) is
        variable readready_v : std_logic;
        begin
            if I_areset = '1' then
                readready_v := '0';
            elsif rising_edge(I_clk) then
                if readready_v = '1' then
                    readready_v := '0';
                elsif I_csboot = '1' then
                    readready_v := '1';
                else
                    readready_v := '0';
                end if;
            end if;

            O_memready <= readready_v;
        end process;
        
    end generate;

    gen_bootrom_not: if not HAVE_BOOTLOADER_ROM generate
        O_load_misaligned_error <= '0';
        O_dataout <= (others => 'X');
        O_instr  <= (others => 'X');
        O_memready <= '0';
    end generate;
end architecture rtl;
