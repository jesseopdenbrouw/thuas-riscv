-- #################################################################################################
-- # io.vhd - The I/O                                                                              #
-- # ********************************************************************************************* #
-- # This file is part of the THUAS RISCV RV32 Project                                             #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2024, Jesse op den Brouw. All rights reserved.                                  #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # https:/github.com/jesseopdenbrouw/thuas-riscv                                                 #
-- #################################################################################################

-- The I/O consists of:
-- A single 32 bits input register and a single 32 bit output
-- register. There is no data direction register. This may be
-- updated in the future. A simple external input interrupt is
-- provided, selecting one of the 32 inputs and rising/falling/both
-- edges.
-- One UART with 7/8/9 data bits, N/E/O parity and 1/2 stop
-- bits. Several UART flags are available: transmit complete,
-- receive complete, parity error, receive failed and framing
-- error. Interrupts on Transmit complete and Receive complete.
-- A simple timer TIMER1 is provided, has no prescaler and
-- generates an interrupt when the CMPT register is equal to
-- or greater than the TCNT register.
-- A more elaborate timer TIMER2 is provided with a 16-bit prescaler
-- PRSC and a 16-bit counter CMPT. Three PWM/OC outputs (A,B,C)
-- are provided. Interrupts available on T/A/B/C.
-- Two minimal I2C master-only devices, I2C1 & I2C2, capable of
-- using Standard mode (Sm) and Fast mode (Fm). START and STOP
-- conditions generated by software settings. Transmit complete
-- interrupt available for I2C1 only.
-- A SPI master device in available, with hardware active low
-- slave select, transmitting 8/16/24/32 bits in one transmission
-- and has interrupt capabilities.
-- A second simple SPI master is included without hardware slave
-- select and no interrupt capabilities.
-- The TIME and TIMECMP registers are provided and are memory
-- mapped and available as output. The TIME registers are currently
-- not writable. 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.processor_common.all;

entity io is
    generic (
          -- The frequency of the system
          SYSTEM_FREQUENCY : integer;
          -- Frequency of the clock (1 MHz)_
          CLOCK_FREQUENCY : integer;
          -- Do we use fast store?
          HAVE_FAST_STORE : boolean;
          -- Do we have UART1?
          HAVE_UART1 : boolean;
          -- Do we have SPI1?
          HAVE_SPI1 : boolean;
          -- Do we have SPI2?
          HAVE_SPI2 : boolean;
          -- Do we have I2C1?
          HAVE_I2C1 : boolean;
          -- Do we have I2C2?
          HAVE_I2C2 : boolean;
          -- Do we have TIMER1?
          HAVE_TIMER1 : boolean;
          -- Do we have TIMER2?
          HAVE_TIMER2 : boolean
         );             
    port (I_clk : in std_logic;
          I_areset : in std_logic;
          I_memaddress : in data_type;
          I_memsize : memsize_type;
          I_csio : in std_logic;
          I_wren : in std_logic;
          I_datain : in data_type;
          O_dataout : out data_type;
          O_memready : out std_logic;
          -- Misaligned access
          O_load_misaligned_error : out std_logic;
          O_store_misaligned_error : out std_logic;
          -- Connection with outside world
          -- GPIOA
          I_gpioapin : in data_type;
          O_gpioapout : out data_type;
          -- UART1
          I_uart1rxd : in std_logic;
          O_uart1txd : out std_logic;
          -- I2C1
          IO_i2c1scl : inout std_logic;
          IO_i2c1sda : inout std_logic;
          -- I2C2
          IO_i2c2scl : inout std_logic;
          IO_i2c2sda : inout std_logic;
          -- SPI1
          O_spi1sck : out std_logic;
          O_spi1mosi : out std_logic;
          I_spi1miso : in std_logic;
          O_spi1nss : out std_logic;
          -- SPI2
          O_spi2sck : out std_logic;
          O_spi2mosi : out std_logic;
          I_spi2miso : in std_logic;
          -- TIMER2
          O_timer2oct : out std_logic;
          IO_timer2icoca : inout std_logic;
          IO_timer2icocb : inout std_logic;
          IO_timer2icocc : inout std_logic;
          -- TIME and TIMEH
          O_mtime : out data_type;
          O_mtimeh : out data_type;
          -- Hardware interrupt request
          O_intrio : out data_type
         );
end entity io;
    
architecture rtl of io is

-- The I/O
-- NOTE: the I/O is word (32 bits) size, Big Endian
--       so there is no need to recode the data
--       The I/O can only handle word size access
--       Set io_size_bits as if it were bytes
-- Default 256 bytes data
constant io_size_bits : integer := 8;
constant io_size : integer := 2**(io_size_bits-2);
type io_type is array (0 to io_size-1) of data_type;

-- The I/O register file, for simulation only
-- synthesis translate_off
signal io_alt : io_type;
-- synthesis translate_on


-- The I/O register number from address
signal reg_int : integer range 0 to io_size-1;
-- Boolean TRUE if the address is on word boundary
signal isword : boolean;
-- Read access granted
signal read_access_granted : std_logic;
-- Write access granted
signal write_access_granted : std_logic;
-- Flop to wait for second read_access_granted (LOAD)
signal read_access_granted_ff : std_logic;
-- Signal is active in second LOAD cycle (read access)
signal read_access_granted_second_cycle : std_logic;
-- Read ready
signal readready : std_logic;

-- Port input and output
constant gpioapin_addr : integer := 0;   -- 0x00.b
constant gpioapout_addr : integer := 1;  -- 0x04.b
constant gpioaextc_addr : integer := 6;  -- 0x18.b
constant gpioaexts_addr : integer := 7;  -- 0x1c.b

type gpioa_type is record
    pin  : data_type;
    pout : data_type;
    extc : data_type;
    exts : data_type;
    pin_sync : data_type;
    ext_sync : std_logic_vector(2 downto 0);
end record;    
signal gpioa : gpioa_type;
-- Note: registers 2 - 5 not used -- reserved


-- UART1
constant uart1ctrl_addr : integer := 8;   -- 0x20.b
constant uart1stat_addr : integer := 9;   -- 0x24.b
constant uart1data_addr : integer := 10;  -- 0x28.b
constant uart1baud_addr : integer := 11;  -- 0x2c.b

type uarttxstate_type is (tx_idle, tx_iter, tx_ready);
type uartrxstate_type is (rx_idle, rx_wait, rx_iter, rx_parity, rx_parity2, rx_ready, rx_fail);

type uart1_type is record
    ctrl : data_type;
    stat : data_type;
    data : data_type;
    baud : data_type;
    -- Transmit signals
    txbuffer : std_logic_vector(11 downto 0);
    txstart : std_logic;
    txstate : uarttxstate_type;
    txbittimer : integer range 0 to 65535;
    txshiftcounter : integer range 0 to 15;
    --Receive signals
    rxbuffer : std_logic_vector(11 downto 0);
    rxstate : uartrxstate_type;
    rxbittimer : integer range 0 to 65535;
    rxshiftcounter : integer range 0 to 15;
    rxd_sync : std_logic;
end record;
signal uart1 : uart1_type;

alias uart1size : std_logic_vector(1 downto 0) is uart1.ctrl(3 downto 2);
alias uart1paron : std_logic is uart1.ctrl(5);
alias uart1parnevenodd : std_logic is uart1.ctrl(4);
alias uart1stop2 : std_logic is uart1.ctrl(0);
alias uart1tc : std_logic is uart1.stat(4);
alias uart1pe : std_logic is uart1.stat(3);
alias uart1rc : std_logic is uart1.stat(2);
alias uart1rf : std_logic is uart1.stat(1);
alias uart1fe : std_logic is uart1.stat(0);

-- Register 12 - 15 not used, reserved


-- I2C1 - minimalistic I2C master-only
constant i2c1ctrl_addr : integer := 16;   -- 0x40.b
constant i2c1stat_addr : integer := 17;   -- 0x44.b
constant i2c1data_addr : integer := 18;   -- 0x48.b

type i2cstate_type is (idle, send_startbit, send_data_first, send_data_second, leadout,
                        send_stopbit_first, send_stopbit_second, send_stopbit_third);
type i2c_type is record
    ctrl : data_type;
    stat : data_type;
    data : data_type;
    state : i2cstate_type;
    bittimer : integer range 0 to 65535;
    shiftcounter : integer range 0 to 9;
    startstransmission : std_logic;
    txbuffer : std_logic_vector(8 downto 0);
    rxbuffer : std_logic_vector(8 downto 0);
    sda_out : std_logic;
    scl_out : std_logic;
    sdasync : std_logic_vector(1 downto 0);
    sclsync : std_logic_vector(1 downto 0);
end record;
signal i2c1 : i2c_type;

alias i2c1mack : std_logic is i2c1.ctrl(11);
alias i2c1hardstop : std_logic is i2c1.ctrl(10);
alias i2c1startbit : std_logic is i2c1.ctrl(9);
alias i2c1stopbit : std_logic is i2c1.ctrl(8);
alias i2c1fastmode : std_logic is i2c1.ctrl(2);
alias i2c1softreset : std_logic is i2c1.ctrl(1);
alias i2c1istransmitting : std_logic is i2c1.stat(2);
alias i2c1tc : std_logic is i2c1.stat(3); 
alias i2c1ackfail : std_logic is i2c1.stat(5);
alias i2c1busy : std_logic is i2c1.stat(6);

-- Register 19 not used, reserved

-- I2C2 - minimalistic I2C master-only
constant i2c2ctrl_addr : integer := 20;   -- 0x50.b
constant i2c2stat_addr : integer := 21;   -- 0x54.b
constant i2c2data_addr : integer := 22;   -- 0x58.b

signal i2c2 : i2c_type;

alias i2c2mack : std_logic is i2c2.ctrl(11);
alias i2c2hardstop : std_logic is i2c2.ctrl(10);
alias i2c2startbit : std_logic is i2c2.ctrl(9);
alias i2c2stopbit : std_logic is i2c2.ctrl(8);
alias i2c2fastmode : std_logic is i2c2.ctrl(2);
alias i2c2softreset : std_logic is i2c2.ctrl(1);
alias i2c2istransmitting : std_logic is i2c2.stat(2);
alias i2c2tc : std_logic is i2c2.stat(3); 
alias i2c2ackfail : std_logic is i2c2.stat(5);
alias i2c2busy : std_logic is i2c2.stat(6);


-- SPI1 - full SPI master with hardware NSS
constant spi1ctrl_addr : integer := 24; -- 0x60.b
constant spi1stat_addr : integer := 25; -- 0x64.b
constant spi1data_addr : integer := 26; -- ox68.b
constant spi1mosidefault : std_logic := 'Z';

type spi1state_type is (idle, cssetup, first, second, leadout, cshold);

type spi1_type is record
    ctrl : data_type;
    stat : data_type;
    data : data_type;
    start : std_logic;
    state : spi1state_type;
    txbuffer : data_type;
    rxbuffer : data_type;
    bittimer : integer range 0 to 127;
    shiftcounter : integer range 0 to 32;
    mosi : std_logic;
    sck : std_logic;
end record;
signal spi1 : spi1_type;
-- Register 27 not used - reserved


-- SPI2 - simple SPI master, software NSS
constant spi2ctrl_addr : integer := 28; -- 0x70.b
constant spi2stat_addr : integer := 29; -- 0x74.b
constant spi2data_addr : integer := 30; -- ox78.b
-- Register 31 not used
constant spi2mosidefault : std_logic := '1';

type spi2state_type is (idle, first, second, leadout);

type spi2_type is record
    ctrl : data_type;
    stat : data_type;
    data : data_type;
    start : std_logic;
    state : spi2state_type;
    txbuffer : data_type;
    rxbuffer : data_type;
    bittimer : integer range 0 to 127;
    shiftcounter : integer range 0 to 32;
    mosi : std_logic;
    sck : std_logic;
end record;
signal spi2 : spi2_type;

-- Register 31 not used - reserved


-- Timer/Counters
-- TIMER1
constant timer1ctrl_addr : integer := 32; -- 0x80.b
constant timer1stat_addr : integer := 33; -- 0x84.b
constant timer1cntr_addr : integer := 34; -- 0x88.b
constant timer1cmpt_addr : integer := 35; -- 0x8c.b
type timer1_type is record
    ctrl : data_type;
    stat : data_type;
    cntr : data_type;
    cmpt : data_type;
end record;
signal timer1 : timer1_type;

-- registers 36 - 39 not used -- reserved


-- TIMER2
constant timer2ctrl_addr : integer := 40; -- 0xa0.b
constant timer2stat_addr : integer := 41; -- 0xa4.b
constant timer2cntr_addr : integer := 42; -- 0xa8.b
constant timer2cmpt_addr : integer := 43; -- 0xac.b
constant timer2prsc_addr : integer := 44; -- 0xb0.b
constant timer2cmpa_addr : integer := 45; -- 0xb4.b
constant timer2cmpb_addr : integer := 46; -- 0xb8.b
constant timer2cmpc_addr : integer := 47; -- 0xbc.b

type timer2_type is record
    ctrl : data_type;
    stat : data_type;
    cntr : data_type;
    cmpt : data_type;
    prsc : data_type;
    cmpa : data_type;
    cmpb : data_type;
    cmpc : data_type;
-- internal prescaler
    prescaler : data_type;
-- shadow registers
    cmptshadow : data_type;
    cmpashadow : data_type;
    cmpbshadow : data_type;
    cmpcshadow : data_type;
    prscshadow : data_type;
    oct : std_logic;
    oca : std_logic;
    ocb : std_logic;
    occ : std_logic;
    ocaen : std_logic;
    ocben : std_logic;
    occen : std_logic;
    icasync : std_logic_vector(2 downto 0);
    icbsync : std_logic_vector(2 downto 0);
    iccsync : std_logic_vector(2 downto 0);
end record;
signal timer2 : timer2_type;

-- Registers 48 - 58 not used - reserved

constant msitrig_addr : integer := 59; -- 0xec.b

-- RISC-V Machine Software Interrupt (MSI)
type msi_type is record
    trig : data_type;
end record;
signal msi : msi_type;

-- RISC-V system timer TIME and TIMECMP
constant mtime_addr : integer := 60;      -- 0xf0.b
constant mtimeh_addr : integer := 61;     -- 0xf4.b
constant mtimecmp_addr : integer := 62;   -- 0xf8.b
constant mtimecmph_addr : integer := 63;  -- 0xfc.b

type mtime_type is record
    mtime : data_type;
    mtimeh : data_type;
    mtimecmp : data_type;
    mtimecmph : data_type;
end record;
signal mtime : mtime_type;

begin

    -- Fetch internal register of io_size_bits bits minus 2
    -- because we will use word size only
    reg_int <= to_integer(unsigned(I_memaddress(io_size_bits-1 downto 2)));
    
    -- Check if an access is on a 4-byte boundary AND is word size
    isword <= TRUE when I_memsize = memsize_word and I_memaddress(1 downto 0) = "00" else FALSE;

    -- Misaligned error, when (not on a 4-byte boundary OR not word size) AND chip select
    O_load_misaligned_error <= '1' when not isword and I_csio = '1' and I_wren = '0' else '0';
    O_store_misaligned_error <= '1' when not isword and I_csio = '1' and I_wren = '1' else '0';
    
    -- Read or write access
    read_access_granted <= '1' when isword and I_csio = '1' and I_wren = '0' else '0';
    write_access_granted <= '1' when isword and I_csio = '1' and I_wren = '1' else '0';
    

    --
    -- Data out to ALU
    --
    process (I_clk, I_areset) is
    begin
        -- Reading a register here doesn't have side effects such as clearing bits.
        if I_areset = '1' then
            O_dataout <= (others => '0');
        elsif rising_edge(I_clk) then
            if read_access_granted = '1' then
                case reg_int is
                    when gpioapin_addr   => O_dataout <= gpioa.pin;
                    when gpioapout_addr  => O_dataout <= gpioa.pout;
                    when gpioaextc_addr  => O_dataout <= gpioa.extc;
                    when gpioaexts_addr  => O_dataout <= gpioa.exts;
                    when uart1ctrl_addr  => O_dataout <= uart1.ctrl;
                    when uart1stat_addr  => O_dataout <= uart1.stat;
                    when uart1data_addr  => O_dataout <= uart1.data;
                    when uart1baud_addr  => O_dataout <= uart1.baud;
                    when i2c1ctrl_addr   => O_dataout <= i2c1.ctrl;
                    when i2c1stat_addr   => O_dataout <= i2c1.stat;
                    when i2c1data_addr   => O_dataout <= i2c1.data;
                    when i2c2ctrl_addr   => O_dataout <= i2c2.ctrl;
                    when i2c2stat_addr   => O_dataout <= i2c2.stat;
                    when i2c2data_addr   => O_dataout <= i2c2.data;
                    when spi1ctrl_addr   => O_dataout <= spi1.ctrl;
                    when spi1stat_addr   => O_dataout <= spi1.stat;
                    when spi1data_addr   => O_dataout <= spi1.data;
                    when spi2ctrl_addr   => O_dataout <= spi2.ctrl;
                    when spi2stat_addr   => O_dataout <= spi2.stat;
                    when spi2data_addr   => O_dataout <= spi2.data;
                    when timer1ctrl_addr => O_dataout <= timer1.ctrl;
                    when timer1stat_addr => O_dataout <= timer1.stat;
                    when timer1cntr_addr => O_dataout <= timer1.cntr;
                    when timer1cmpt_addr => O_dataout <= timer1.cmpt;
                    when timer2ctrl_addr => O_dataout <= timer2.ctrl;
                    when timer2stat_addr => O_dataout <= timer2.stat;
                    when timer2cntr_addr => O_dataout <= timer2.cntr;
                    when timer2cmpt_addr => O_dataout <= timer2.cmpt;
                    when timer2prsc_addr => O_dataout <= timer2.prsc;
                    when timer2cmpa_addr => O_dataout <= timer2.cmpa;
                    when timer2cmpb_addr => O_dataout <= timer2.cmpb;
                    when timer2cmpc_addr => O_dataout <= timer2.cmpc;
                    when msitrig_addr    => O_dataout <= msi.trig;
                    when mtime_addr      => O_dataout <= mtime.mtime;
                    when mtimeh_addr     => O_dataout <= mtime.mtimeh;
                    when mtimecmp_addr   => O_dataout <= mtime.mtimecmp;
                    when mtimecmph_addr  => O_dataout <= mtime.mtimecmph;
                    when others => O_dataout <= (others => '-');
                end case;
            end if;
        end if;
    end process;

    --
    -- GPIO A pin en pout    
    -- General purpose I/O ports, one 32-bit input and one 32-bit output
    --
    process (I_clk, I_areset) is
    begin
        if I_areset = '1' then
            gpioa.pin <= (others => '0');
            gpioa.pout <= (others => '0');
            gpioa.pin_sync <= (others => '0');
            gpioa.extc <= (others => '0');
            gpioa.exts <= (others => '0');
            gpioa.ext_sync <= (others => '0');
        elsif rising_edge(I_clk) then
            -- Read data in from outside world
            -- Synchronizer register
            gpioa.pin_sync <= I_gpioapin; 
            gpioa.pin <= gpioa.pin_sync;
            -- External interrupt
            gpioa.ext_sync <= gpioa.ext_sync(1 downto 0) & I_gpioapin(to_integer(unsigned(gpioa.extc(7 downto 3))));
            -- Only write to I/O when write is enabled AND size is word
            -- Only write to the outputs, not the inputs
            -- Only write if on 4-byte boundary
            -- Only write when Chip Select (cs)
            if write_access_granted = '1' then
                if reg_int = gpioapout_addr then
                    gpioa.pout <= I_datain;
                elsif reg_int = gpioaextc_addr then
                    gpioa.extc <= I_datain;
                elsif reg_int = gpioaexts_addr then
                    gpioa.exts <= I_datain;
                end if;
            end if;
            -- Detect rising edge or falling edge or both
            if (gpioa.extc(1) = '1' and gpioa.ext_sync(2) = '0' and gpioa.ext_sync(1) = '1') or
               (gpioa.extc(2) = '1' and gpioa.ext_sync(2) = '1' and gpioa.ext_sync(1) = '0') then
                gpioa.exts(0) <= '1';
            end if;
        end if;
    end process;
     -- Data to outside world
    O_gpioapout <= gpioa.pout;
    
    
    --
    -- UART1
    --
    uart1gen: if HAVE_UART1 generate
        process (I_clk, I_areset) is
        variable uart1txshiftcounter_var : integer range 0 to 15;
        begin
            -- Common resets et al.
            if I_areset = '1' then
                uart1.data <= (others => '0');
                uart1.baud <= (others => '0');
                uart1.ctrl <= (others => '0');
                uart1.stat <= (others => '0');
                uart1.txstart <= '0';
                uart1.txstate <= tx_idle;
                uart1.txbuffer <= (others => '0');
                uart1.txbittimer <= 0;
                uart1.txshiftcounter <= 0;
                O_uart1txd <= '1';
                uart1.rxbuffer <= (others => '0');
                uart1.rxstate <= rx_idle;
                uart1.rxbittimer <= 0;
                uart1.rxshiftcounter <= 0;
                uart1.rxd_sync <= '1';
            elsif rising_edge(I_clk) then
                -- Default for start transmission
                uart1.txstart <= '0';
                -- Common register writes
                if write_access_granted = '1' then
                    if reg_int = uart1ctrl_addr then
                        -- A write to the control register
                        uart1.ctrl <= I_datain;
                    elsif reg_int = uart1stat_addr then
                        -- A write to the status register
                        uart1.stat <= I_datain;
                    elsif reg_int = uart1baud_addr then
                        -- A write to the baud rate register
                        -- Use only 16 bits for baud rate
                        uart1.baud <= I_datain;
                    elsif reg_int = uart1data_addr then
                        -- A write to the data register triggers a transmission
                        -- Signal start
                        uart1.txstart <= '1';
                        -- Load transmit buffer with 7/8/9 data bits, parity bit and
                        -- a start bit
                        -- Stop bits will be automatically added since the remaining
                        -- bits are set to 1. Most right bit is start bit.
                        uart1.txbuffer <= (others => '1');
                        if uart1size = "10" then
                            -- 9 bits data
                            uart1.txbuffer(9 downto 0) <= I_datain(8 downto 0) & '0';
                            -- Have parity
                            if uart1paron = '1' then
                                uart1.txbuffer(10) <= I_datain(8) xor I_datain(7) xor I_datain(6) xor I_datain(5) xor I_datain(4)
                                                  xor I_datain(3) xor I_datain(2) xor I_datain(1) xor I_datain(0) xor uart1parnevenodd;
                            end if;
                        elsif uart1size = "11" then
                            -- 7 bits data
                            uart1.txbuffer(7 downto 0) <= I_datain(6 downto 0) & '0';
                            -- Have parity
                            if uart1paron = '1' then
                                uart1.txbuffer(8) <= I_datain(6) xor I_datain(5) xor I_datain(4) xor I_datain(3)
                                                 xor I_datain(2) xor I_datain(1) xor I_datain(0) xor uart1parnevenodd;
                            end if;
                        else
                            -- 8 bits data
                            uart1.txbuffer(8 downto 0) <= I_datain(7 downto 0) & '0';
                            -- Have parity
                            if uart1paron = '1' then
                                uart1.txbuffer(9) <= I_datain(7) xor I_datain(6) xor I_datain(5) xor I_datain(4) xor I_datain(3)
                                                 xor I_datain(2) xor I_datain(1) xor I_datain(0) xor uart1parnevenodd;
                            end if;
                        end if;
                        -- Signal that we are sending
                        uart1tc <= '0'; 
                    end if;
                end if;
                
                -- If data register is read...
                -- Reading data register clears flags!
                if read_access_granted_second_cycle = '1' then
                    if reg_int = uart1data_addr then
                        -- Clear the received status bits
                        -- PE, RC, RF, FE
                        uart1pe <= '0';
                        uart1rc <= '0';
                        uart1rf <= '0';
                        uart1fe <= '0';
                    end if;
                end if;
                
                -- Transmit a character
                case uart1.txstate is
                    -- Tx idle state, wait for start
                    when tx_idle =>
                        O_uart1txd <= '1';
                        -- If start triggered...
                        if uart1.txstart = '1' then
                            -- Load the prescaler, set the number of bits (including start bit)
                            uart1.txbittimer <= to_integer(unsigned(uart1.baud));
                            if uart1size = "10" then
                                uart1txshiftcounter_var := 10;
                            elsif uart1size = "11" then
                                uart1txshiftcounter_var := 8;
                            else
                                uart1txshiftcounter_var := 9;
                            end if;
                            -- Add up possible parity bit and possible second stop bit
                            if uart1paron = '1' then
                                uart1txshiftcounter_var := uart1txshiftcounter_var + 1;
                            end if;
                            if uart1stop2 = '1' then
                                uart1txshiftcounter_var := uart1txshiftcounter_var + 1;
                            end if;
                            uart1.txshiftcounter <= uart1txshiftcounter_var;
                            uart1.txstate <= tx_iter;
                        else
                            uart1.txstate <= tx_idle;
                        end if;
                    -- Transmit the bits
                    when tx_iter =>
                        -- Cycle through all bits in the transmit buffer
                        -- First in line is the start bit
                        O_uart1txd <= uart1.txbuffer(0);
                        if uart1.txbittimer > 0 then
                            uart1.txbittimer <= uart1.txbittimer - 1;
                        elsif uart1.txshiftcounter > 0 then
                            uart1.txbittimer <= to_integer(unsigned(uart1.baud));
                            uart1.txshiftcounter <= uart1.txshiftcounter - 1;
                            -- Shift in stop bit
                            uart1.txbuffer <= '1' & uart1.txbuffer(uart1.txbuffer'high downto 1);
                        else
                            uart1.txstate <= tx_ready;
                        end if;
                    -- Signal ready
                    when tx_ready =>
                        O_uart1txd <= '1';
                        uart1.txstate <= tx_idle;
                        -- Signal character transmitted
                        uart1tc <= '1'; 
                    when others =>
                        O_uart1txd <= '1';
                        uart1.txstate <= tx_idle;
                end case;
                
                -- Receive character
                -- Input synchronizer
                uart1.rxd_sync <= I_uart1rxd;
                case uart1.rxstate is
                    -- Rx idle, wait for start bit
                    when rx_idle =>
                        -- If detected a start bit ...
                        if uart1.rxd_sync = '0' then
                            -- Set half bit time ...
                            uart1.rxbittimer <= to_integer(unsigned(uart1.baud))/2;
                            uart1.rxstate <= rx_wait;
                        else
                            uart1.rxstate <= rx_idle;
                        end if;
                    -- Hunt for start bit, check start bit at half bit time
                    when rx_wait =>
                        if uart1.rxbittimer > 0 then
                            uart1.rxbittimer <= uart1.rxbittimer - 1;
                        else
                            -- At half bit time...
                            -- Start bit is still 0, so continue
                            if uart1.rxd_sync = '0' then
                                uart1.rxbittimer <= to_integer(unsigned(uart1.baud));
                                -- Set reception size
                                if uart1size = "10" then
                                    -- 9 bits
                                    uart1.rxshiftcounter <= 9;
                                elsif uart1size = "11" then
                                    -- 7 bits
                                    uart1.rxshiftcounter <= 7;
                                else
                                    -- 8 bits
                                    uart1.rxshiftcounter <= 8;
                                end if;
                                uart1.rxbuffer <= (others => '0');
                                uart1.rxstate <= rx_iter;
                            else
                                -- Start bit is not 0, so invalid transmission
                                uart1.rxstate <= rx_fail;
                            end if;
                        end if;
                    -- Shift in the data bits
                    -- We sample in the middle of a bit time...
                    when rx_iter =>
                        if uart1.rxbittimer > 0 then
                            -- Bit timer not finished, so keep counting...
                            uart1.rxbittimer <= uart1.rxbittimer - 1;
                        elsif uart1.rxshiftcounter > 0 then
                            -- Bit counter not finished, so restart timer and shift in data bit
                            uart1.rxbittimer <= to_integer(unsigned(uart1.baud));
                            uart1.rxshiftcounter <= uart1.rxshiftcounter - 1;
                            if uart1size = "10" then
                                -- 9 bits
                                uart1.rxbuffer(8 downto 0) <= uart1.rxd_sync & uart1.rxbuffer(8 downto 1);
                            elsif uart1size = "11" then
                                -- 7 bits
                                uart1.rxbuffer(6 downto 0) <= uart1.rxd_sync & uart1.rxbuffer(6 downto 1);
                            else
                                -- 8 bits
                                uart1.rxbuffer(7 downto 0) <= uart1.rxd_sync & uart1.rxbuffer(7 downto 1);
                            end if;
                        else
                            -- Do we have a parity bit?
                            if uart1paron = '1' then
                                uart1.rxstate <= rx_parity;
                            else
                                uart1.rxstate <= rx_ready;
                            end if;
                        end if;
                    -- Check parity, we already there...
                    when rx_parity =>
                        if uart1size = "10" then
                            uart1pe <= uart1.rxbuffer(8) xor uart1.rxbuffer(7) xor uart1.rxbuffer(6) xor uart1.rxbuffer(5)
                                                xor uart1.rxbuffer(4) xor uart1.rxbuffer(3) xor uart1.rxbuffer(2)
                                                xor uart1.rxbuffer(1) xor uart1.rxbuffer(0) xor uart1.rxd_sync xor uart1parnevenodd;
                        elsif uart1size = "11" then
                            uart1pe <= uart1.rxbuffer(6) xor uart1.rxbuffer(5)
                                                xor uart1.rxbuffer(4) xor uart1.rxbuffer(3) xor uart1.rxbuffer(2)
                                                xor uart1.rxbuffer(1) xor uart1.rxbuffer(0) xor uart1.rxd_sync xor uart1parnevenodd;
                        else
                            uart1pe <= uart1.rxbuffer(7) xor uart1.rxbuffer(6) xor uart1.rxbuffer(5)
                                                xor uart1.rxbuffer(4) xor uart1.rxbuffer(3) xor uart1.rxbuffer(2)
                                                xor uart1.rxbuffer(1) xor uart1.rxbuffer(0) xor uart1.rxd_sync xor uart1parnevenodd;
                        end if;
                        uart1.rxbittimer <= to_integer(unsigned(uart1.baud));
                        uart1.rxstate <= rx_parity2;
                    -- Wait to middle of stop bit
                    when rx_parity2 =>
                        if uart1.rxbittimer > 0 then
                            uart1.rxbittimer <= uart1.rxbittimer - 1;
                        else
                            uart1.rxstate <= rx_ready;
                        end if;
                    -- When ready, all bits are shifted in
                    -- Even if we use two stop bits, we only check one and
                    -- signal reception. This leave some computation time
                    -- before the next reception occurs.
                    when rx_ready =>
                        -- Test for a stray 0 in position of (first) stop bit
                        if uart1.rxd_sync = '0' then
                            -- Signal frame error
                            uart1fe <= '1';
                        end if;
                        -- Any way, copy the received data to the data register
                        uart1.data <= (others => '0');
                        if uart1size = "10" then
                            -- 9 bits
                            uart1.data(8 downto 0) <= uart1.rxbuffer(8 downto 0);
                        elsif uart1size = "11" then
                            -- 7 bits
                            uart1.data(6 downto 0) <= uart1.rxbuffer(6 downto 0);
                        else
                            -- 8 bits
                            uart1.data(7 downto 0) <= uart1.rxbuffer(7 downto 0);
                        end if;
                        -- signal reception
                        uart1rc <= '1';
                        uart1.rxstate <= rx_idle;
                    -- Wrong start bit detected, no data present
                    when rx_fail =>
                        -- Failed to receive a correct start bit...
                        uart1.rxstate <= rx_idle;
                        uart1rf <= '1';
                    when others =>
                        uart1.rxstate <= rx_idle;
                end case;
                uart1.baud(31 downto 16) <= (others => '0');
                uart1.data(31 downto 9) <= (others => '0');
                uart1.ctrl(31 downto 8) <= (others => '0');
                uart1.stat(31 downto 5) <= (others => '0');
            end if;
        end process;
    end generate;
    uart1gen_not: if not HAVE_UART1 generate
        uart1.baud <= (others => '0');
        uart1.data <= (others => '0');
        uart1.ctrl <= (others => '0');
        uart1.stat <= (others => '0');
        O_uart1txd <= 'Z';
    end generate;

    --
    -- I2C1
    --
    i2c1gen : if HAVE_I2C1 generate
        process (I_clk, I_areset) is
        begin
            if I_areset = '1' then
                i2c1.ctrl <= (others => '0');
                i2c1.stat <= (others => '0');
                i2c1.data <= (others => '0');
                i2c1.scl_out <= '1';
                i2c1.sda_out <= '1';
                i2c1.state <= idle;
                i2c1.bittimer <= 0;
                i2c1.shiftcounter <= 0;
                i2c1.txbuffer <= (others => '0');
                i2c1.rxbuffer <= (others => '0');
                i2c1.startstransmission <= '0';
                i2c1.sclsync <= (others => '1');
                i2c1.sdasync <= (others => '1');
            elsif rising_edge(I_clk) then
                i2c1.startstransmission <= '0';
                -- Common register writes
                if write_access_granted = '1' then
                    if reg_int = i2c1ctrl_addr then
                        i2c1.ctrl <= I_datain;
                    elsif reg_int = i2c1stat_addr then
                        i2c1.stat <= I_datain;
                    elsif reg_int = i2c1data_addr then
                        -- Latch data, if startbit set, end with master Nack
                        i2c1.txbuffer <= I_datain(7 downto 0) & (i2c1startbit or i2c1stopbit or not i2c1mack);
                        -- Signal that we are sending data
                        i2c1.startstransmission <= '1';
                        -- Reset both Transmission Complete and Ack Failed
                        i2c1tc <= '0';
                        i2c1ackfail <= '0';
                    end if;
                end if;
                -- If read data register, clear the TC and AF flag
                -- Reading data register clears flags!
                if read_access_granted_second_cycle = '1' then
                    if reg_int = i2c1data_addr then
                        i2c1tc <= '0';
                        i2c1ackfail <= '0';
                    end if;
                end if;

                -- Check for I2C bus is busy.
                -- If SCL or SDA is/are low...
                if i2c1.sclsync(1) = '0' or i2c1.sdasync(1) = '0' then
                    -- I2C bus is busy
                    i2c1busy <= '1';
                end if;
                -- SCL is high and rising edge on SDA...
                if i2c1.sclsync(0) /= '0' and i2c1.sdasync(1) = '0' and i2c1.sdasync(0) /= '0' then
                    -- signals a STOP, so bus is free
                    i2c1busy <= '0';
                end if;
                
                -- Input synchronizer
                i2c1.sdasync <= i2c1.sdasync(0) & IO_i2c1sda;
                i2c1.sclsync <= i2c1.sclsync(0) & IO_i2c1scl;

                -- The I2C1 state machine
                case i2c1.state is
                    when idle =>
                        -- Clock == !state_of_transmitting, SDA = High-Z (==1)
                        -- If transmitting, the clock is held low. If not
                        -- transmitting, the clock is held high (high-Z). After
                        -- STOP, the state of transmitting is reset. This keeps
                        -- the bus occupied between START and STOP.
                        i2c1.scl_out <= not i2c1istransmitting;
                        i2c1.sda_out <= '1';
                        -- Idle situation, load the counters and set SCL/SDA to High-Z
                        if i2c1fastmode = '1' then
                            i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)))*2;
                        else
                            i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)));
                        end if;
                        i2c1.shiftcounter <= 8;
                        -- Is data register written?
                        if i2c1.startstransmission = '1' then
                            -- Register that we are transmitting
                            i2c1istransmitting <= '1';
                            -- Data written to data register, check for start condition
                            if i2c1startbit = '1' then
                                -- Start bit is seen, so clear it.
                                i2c1startbit <= '0';
                                -- Send a START bit, so address comes next
                                i2c1.state <= send_startbit;
                            else
                                -- Regular data
                                i2c1.state <= send_data_first;
                            end if;
                        -- Do we have to send a single STOP condition?
                        elsif i2c1hardstop = '1' then
                            i2c1.state <= send_stopbit_first;
                        end if;
                    when send_startbit =>
                        -- Generate start condition
                        i2c1.scl_out <= '1';
                        i2c1.sda_out <= '0';
                        if i2c1.bittimer > 0 then
                            i2c1.bittimer <= i2c1.bittimer - 1;
                        else
                            if i2c1fastmode = '1' then
                                i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)))*2;
                            else
                                i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)));
                            end if;
                            i2c1.state <= send_data_first;
                        end if;
                    when send_data_first =>
                        -- SCL low == 0, SDA 0 or High-Z (== 1)
                        i2c1.scl_out <= '0';
                        i2c1.sda_out <= i2c1.txbuffer(8);
                        
                        -- Count bit time
                        if i2c1.bittimer > 0 then
                            i2c1.bittimer <= i2c1.bittimer - 1;
                        else
                            i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)));
                            i2c1.state <= send_data_second;
                        end if;
                    when send_data_second =>
                        -- SCL High-Z == 1, SDA 0 or High-Z (== 1)
                        i2c1.scl_out <= '1';
                        i2c1.sda_out <= i2c1.txbuffer(8);

                        -- Count bit time
                        if i2c1.bittimer > 0 then
                            i2c1.bittimer <= i2c1.bittimer - 1;
                        else
                            if i2c1fastmode = '1' then
                                i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)))*2;
                            else
                                i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)));
                            end if;
                            -- Check if more bits
                            if i2c1.shiftcounter > 0 then
                                -- More bits to send...
                                i2c1.shiftcounter <= i2c1.shiftcounter - 1;
                                i2c1.state <= send_data_first;
                                -- Shift next bit, hold time is 0 ns as per spec
                                i2c1.txbuffer <= i2c1.txbuffer(7 downto 0) & '1';
                            else
                                -- No more bits, then goto STOP or leadout
                                if i2c1stopbit = '1' then
                                    i2c1.state <= send_stopbit_first;
                                else
                                    i2c1.state <= leadout;
                                end if;
                            end if;
                        end if;
                        -- If detected rising edge on external SCL, clock in SDA.
                        if i2c1.sclsync(1) = '0' and i2c1.sclsync(0) /= '0' then
                            i2c1.rxbuffer <= i2c1.rxbuffer(7 downto 0) & i2c1.sdasync(1);
                        end if;
                    when leadout =>
                        -- SCL low, SDA high
                        i2c1.scl_out <= '0';
                        i2c1.sda_out <= '1';
                        -- Count bit time
                        if i2c1.bittimer > 0 then
                            i2c1.bittimer <= i2c1.bittimer - 1;
                        else
                            --i2c1bittimer <= to_integer(unsigned(i2c1ctrl_int(31 downto 16)));
                            i2c1.state <= idle;
                            i2c1tc <= '1';
                            i2c1.data(7 downto 0) <= i2c1.rxbuffer(8 downto 1);
                            i2c1ackfail <= i2c1.rxbuffer(0);
                        end if;
                    when send_stopbit_first =>
                        -- SCL low, SDA low
                        i2c1.scl_out <= '0';
                        i2c1.sda_out <= '0';
                        -- Count bit time
                        if i2c1.bittimer > 0 then
                            i2c1.bittimer <= i2c1.bittimer - 1;
                        else
                            i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)));
                            i2c1.state <= send_stopbit_second;
                        end if;
                    when send_stopbit_second =>
                        -- SCL high, SDA low
                        i2c1.scl_out <= '1';
                        i2c1.sda_out <= '0';
                        -- Count bit timer
                        if i2c1.bittimer > 0 then
                            i2c1.bittimer <= i2c1.bittimer - 1;
                        else
                            if i2c1fastmode = '1' then
                                i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)))*2;
                            else
                                i2c1.bittimer <= to_integer(unsigned(i2c1.ctrl(31 downto 16)));
                            end if;
                            i2c1.state <= send_stopbit_third;
                        end if;
                    when send_stopbit_third =>
                        -- SCL high, SCL low, will be set high in idle,
                        -- so there is no need to set SDA high here.
                        i2c1.scl_out <= '1';
                        i2c1.sda_out <= '1';
                        -- Count bit timer
                        if i2c1.bittimer > 0 then
                            i2c1.bittimer <= i2c1.bittimer - 1;
                        else
                            -- Transmission conplete
                            i2c1tc <= '1';
                            -- Clear STOP bit
                            i2c1stopbit <= '0';
                            -- and goto IDLE
                            i2c1.state <= idle;
                            -- Copy data to data register and flag ACK
                            i2c1.data(7 downto 0) <= i2c1.rxbuffer(8 downto 1);
                            i2c1ackfail <= i2c1.rxbuffer(0);
                            -- Clear hard stop
                            i2c1hardstop <= '0';
                            -- Unregister that we are transmitting
                            i2c1istransmitting <= '0';
                        end if;
                    when others =>
                        i2c1.state <= idle;
                end case;
                -- Clear unusd bits
                i2c1.data(31 downto 8) <= (others => '0');
                i2c1.ctrl(15 downto 12) <= (others => '0');
                i2c1.ctrl(7 downto 4) <= (others => '0');
                i2c1.stat(31 downto 12) <= (others => '0');
            end if;
        end process;
        -- Drive the clock and data lines
        IO_i2c1scl <= '0' when i2c1.scl_out = '0' else 'Z';
        IO_i2c1sda <= '0' when i2c1.sda_out = '0' else 'Z';
    end generate;
    i2c1gen_not : if not HAVE_I2C1 generate
        i2c1.data <= (others => '0');
        i2c1.ctrl <= (others => '0');
        i2c1.stat <= (others => '0');
        IO_i2c1scl <= 'Z';
        IO_i2c1sda <= 'Z';
    end generate;

    --
    -- I2C2
    --
    i2c2gen : if HAVE_I2C2 generate
        process (I_clk, I_areset) is
        begin
            if I_areset = '1' then
                i2c2.ctrl <= (others => '0');
                i2c2.stat <= (others => '0');
                i2c2.data <= (others => '0');
                i2c2.scl_out <= '1';
                i2c2.sda_out <= '1';
                i2c2.state <= idle;
                i2c2.bittimer <= 0;
                i2c2.shiftcounter <= 0;
                i2c2.txbuffer <= (others => '0');
                i2c2.rxbuffer <= (others => '0');
                i2c2.startstransmission <= '0';
                i2c2.sclsync <= (others => '1');
                i2c2.sdasync <= (others => '1');
            elsif rising_edge(I_clk) then
                i2c2.startstransmission <= '0';
                -- Common register writes
                if write_access_granted = '1' then
                    if reg_int = i2c2ctrl_addr then
                        i2c2.ctrl <= I_datain;
                    elsif reg_int = i2c2stat_addr then
                        i2c2.stat <= I_datain;
                    elsif reg_int = i2c2data_addr then
                        -- Latch data, if startbit set, end with master Nack
                        i2c2.txbuffer <= I_datain(7 downto 0) & (i2c2startbit or i2c2stopbit or not i2c2mack);
                        -- Signal that we are sending data
                        i2c2.startstransmission <= '1';
                        -- Reset both Transmission Complete and Ack Failed
                        i2c2tc <= '0';
                        i2c2ackfail <= '0';
                    end if;
                end if;
                -- If read data register, clear the TC and AF flag
                -- Reading data register clears flags!
                if read_access_granted_second_cycle = '1' then
                    if reg_int = i2c2data_addr then
                        i2c2tc <= '0';
                        i2c2ackfail <= '0';
                    end if;
                end if;

                -- Check for I2C bus is busy.
                -- If SCL or SDA is/are low...
                if i2c2.sclsync(1) = '0' or i2c2.sdasync(1) = '0' then
                    -- I2C bus is busy
                    i2c2busy <= '1';
                end if;
                -- SCL is high and rising edge on SDA...
                if i2c2.sclsync(0) /= '0' and i2c2.sdasync(1) = '0' and i2c2.sdasync(0) /= '0' then
                    -- signals a STOP, so bus is free
                    i2c2busy <= '0';
                end if;
                
                -- Input synchronizer
                i2c2.sdasync <= i2c2.sdasync(0) & IO_i2c2sda;
                i2c2.sclsync <= i2c2.sclsync(0) & IO_i2c2scl;

                -- The i2c2 state machine
                case i2c2.state is
                    when idle =>
                        -- Clock == !state_of_transmitting, SDA = High-Z (==1)
                        -- If transmitting, the clock is held low. If not
                        -- transmitting, the clock is held high (high-Z). After
                        -- STOP, the state of transmitting is reset. This keeps
                        -- the bus occupied between START and STOP.
                        i2c2.scl_out <= not i2c2istransmitting;
                        i2c2.sda_out <= '1';
                        -- Idle situation, load the counters and set SCL/SDA to High-Z
                        if i2c2fastmode = '1' then
                            i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)))*2;
                        else
                            i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)));
                        end if;
                        i2c2.shiftcounter <= 8;
                        -- Is data register written?
                        if i2c2.startstransmission = '1' then
                            -- Register that we are transmitting
                            i2c2istransmitting <= '1';
                            -- Data written to data register, check for start condition
                            if i2c2startbit = '1' then
                                -- Start bit is seen, so clear it.
                                i2c2startbit <= '0';
                                -- Send a START bit, so address comes next
                                i2c2.state <= send_startbit;
                            else
                                -- Regular data
                                i2c2.state <= send_data_first;
                            end if;
                        -- Do we have to send a single STOP condition?
                        elsif i2c2hardstop = '1' then
                            i2c2.state <= send_stopbit_first;
                        end if;
                    when send_startbit =>
                        -- Generate start condition
                        i2c2.scl_out <= '1';
                        i2c2.sda_out <= '0';
                        if i2c2.bittimer > 0 then
                            i2c2.bittimer <= i2c2.bittimer - 1;
                        else
                            if i2c2fastmode = '1' then
                                i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)))*2;
                            else
                                i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)));
                            end if;
                            i2c2.state <= send_data_first;
                        end if;
                    when send_data_first =>
                        -- SCL low == 0, SDA 0 or High-Z (== 1)
                        i2c2.scl_out <= '0';
                        i2c2.sda_out <= i2c2.txbuffer(8);
                        
                        -- Count bit time
                        if i2c2.bittimer > 0 then
                            i2c2.bittimer <= i2c2.bittimer - 1;
                        else
                            i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)));
                            i2c2.state <= send_data_second;
                        end if;
                    when send_data_second =>
                        -- SCL High-Z == 1, SDA 0 or High-Z (== 1)
                        i2c2.scl_out <= '1';
                        i2c2.sda_out <= i2c2.txbuffer(8);

                        -- Count bit time
                        if i2c2.bittimer > 0 then
                            i2c2.bittimer <= i2c2.bittimer - 1;
                        else
                            if i2c2fastmode = '1' then
                                i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)))*2;
                            else
                                i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)));
                            end if;
                            -- Check if more bits
                            if i2c2.shiftcounter > 0 then
                                -- More bits to send...
                                i2c2.shiftcounter <= i2c2.shiftcounter - 1;
                                i2c2.state <= send_data_first;
                                -- Shift next bit, hold time is 0 ns as per spec
                                i2c2.txbuffer <= i2c2.txbuffer(7 downto 0) & '1';
                            else
                                -- No more bits, then goto STOP or leadout
                                if i2c2stopbit = '1' then
                                    i2c2.state <= send_stopbit_first;
                                else
                                    i2c2.state <= leadout;
                                end if;
                            end if;
                        end if;
                        -- If detected rising edge on external SCL, clock in SDA.
                        if i2c2.sclsync(1) = '0' and i2c2.sclsync(0) /= '0' then
                            i2c2.rxbuffer <= i2c2.rxbuffer(7 downto 0) & i2c2.sdasync(1);
                        end if;
                    when leadout =>
                        -- SCL low, SDA high
                        i2c2.scl_out <= '0';
                        i2c2.sda_out <= '1';
                        -- Count bit time
                        if i2c2.bittimer > 0 then
                            i2c2.bittimer <= i2c2.bittimer - 1;
                        else
                            --i2c2bittimer <= to_integer(unsigned(i2c2ctrl_int(31 downto 16)));
                            i2c2.state <= idle;
                            i2c2tc <= '1';
                            i2c2.data(7 downto 0) <= i2c2.rxbuffer(8 downto 1);
                            i2c2ackfail <= i2c2.rxbuffer(0);
                        end if;
                    when send_stopbit_first =>
                        -- SCL low, SDA low
                        i2c2.scl_out <= '0';
                        i2c2.sda_out <= '0';
                        -- Count bit time
                        if i2c2.bittimer > 0 then
                            i2c2.bittimer <= i2c2.bittimer - 1;
                        else
                            i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)));
                            i2c2.state <= send_stopbit_second;
                        end if;
                    when send_stopbit_second =>
                        -- SCL high, SDA low
                        i2c2.scl_out <= '1';
                        i2c2.sda_out <= '0';
                        -- Count bit timer
                        if i2c2.bittimer > 0 then
                            i2c2.bittimer <= i2c2.bittimer - 1;
                        else
                            if i2c2fastmode = '1' then
                                i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)))*2;
                            else
                                i2c2.bittimer <= to_integer(unsigned(i2c2.ctrl(31 downto 16)));
                            end if;
                            i2c2.state <= send_stopbit_third;
                        end if;
                    when send_stopbit_third =>
                        -- SCL high, SCL low, will be set high in idle,
                        -- so there is no need to set SDA high here.
                        i2c2.scl_out <= '1';
                        i2c2.sda_out <= '1';
                        -- Count bit timer
                        if i2c2.bittimer > 0 then
                            i2c2.bittimer <= i2c2.bittimer - 1;
                        else
                            -- Transmission conplete
                            i2c2tc <= '1';
                            -- Clear STOP bit
                            i2c2stopbit <= '0';
                            -- and goto IDLE
                            i2c2.state <= idle;
                            -- Copy data to data register and flag ACK
                            i2c2.data(7 downto 0) <= i2c2.rxbuffer(8 downto 1);
                            i2c2ackfail <= i2c2.rxbuffer(0);
                            -- Clear hard stop
                            i2c2hardstop <= '0';
                            -- Unregister that we are transmitting
                            i2c2istransmitting <= '0';
                        end if;
                    when others =>
                        i2c2.state <= idle;
                end case;
                -- Clear unusd bits
                i2c2.data(31 downto 8) <= (others => '0');
                i2c2.ctrl(15 downto 12) <= (others => '0');
                i2c2.ctrl(7 downto 4) <= (others => '0');
                i2c2.stat(31 downto 12) <= (others => '0');
            end if;
        end process;
        -- Drive the clock and data lines
        IO_i2c2scl <= '0' when i2c2.scl_out = '0' else 'Z';
        IO_i2c2sda <= '0' when i2c2.sda_out = '0' else 'Z';
    end generate;
    i2c2gen_not : if not HAVE_I2C2 generate
        i2c2.data <= (others => '0');
        i2c2.ctrl <= (others => '0');
        i2c2.stat <= (others => '0');
        IO_i2c2scl <= 'Z';
        IO_i2c2sda <= 'Z';
    end generate;

    --
    -- SPI1
    --
    spi1gen : if HAVE_SPI1 generate
        process (I_clk, I_areset) is
        variable spi1txshiftcounter_var : integer range 0 to 31;
        variable spi1prescaler_var : integer range 0 to 255;
        begin
            -- Common resets et al.
            if I_areset = '1' then
                spi1.data <= (others => '0');
                spi1.ctrl <= (others => '0');
                spi1.stat <= (others => '0');
                spi1.start <= '0';
                spi1.state <= idle;
                spi1.txbuffer <= (others => '0');
                spi1.bittimer <= 0;
                spi1.shiftcounter <= 0;
                spi1.mosi <= spi1mosidefault;
                spi1.rxbuffer <= (others => '0');
                --spi1miso_sync <= '0';
                spi1.sck <= '0';
                O_spi1nss <= '1';
            elsif rising_edge(I_clk) then
                -- Default for start transmission
                spi1.start <= '0';
                -- Common register writes
                if write_access_granted = '1' then
                    if reg_int = spi1ctrl_addr then
                        -- A write to the control register
                        spi1.ctrl <= I_datain;
                        -- Set clock polarity
                        spi1.sck <= I_datain(2);
                    elsif reg_int = spi1stat_addr then
                        -- A write to the status register
                        spi1.stat <= I_datain;
                    elsif reg_int = spi1data_addr then
                        -- A write to the data register triggers a transmission
                        -- Signal start
                        spi1.start <= '1';
                        -- Load transmit buffer with 8/16/24/32 data bits
                        spi1.txbuffer <= (others => '0');
                        spi1.data <= (others => '0');
                        -- Load the desired bits to transfer
                        case spi1.ctrl(5 downto 4) is
                            when "00" =>   spi1.txbuffer(31 downto 24) <= I_datain(7 downto 0);
                                           spi1.shiftcounter <= 7;
                            when "01" =>   spi1.txbuffer(31 downto 16) <= I_datain(15 downto 0);
                                           spi1.shiftcounter <= 15;
                            when "10" =>   spi1.txbuffer(31 downto 8) <= I_datain(23 downto 0);
                                           spi1.shiftcounter <= 23;
                            when "11" =>   spi1.txbuffer <= I_datain;
                                           spi1.shiftcounter <= 31;
                            when others => spi1.txbuffer <= (others => '-');
                                           spi1.shiftcounter <= 0;
                        end case;
                        -- Signal that we are sending
                        spi1.stat(3) <= '0'; 
                    end if;
                end if;
                -- Zero out bits not needed
                spi1.ctrl(31 downto 28) <= (others => '0');
                spi1.ctrl(11) <= '0';
                spi1.ctrl(7 downto 6) <= (others => '0');
                spi1.ctrl(0) <= '0';
                spi1.stat(31 downto 4) <= (others => '0');
                spi1.stat(2 downto 0) <= (others =>'0');

                -- Calculate prescaler
                case spi1.ctrl(10 downto 8) is
                    when "000" => spi1prescaler_var := 0;
                    when "001" => spi1prescaler_var := 1;
                    when "010" => spi1prescaler_var := 3;
                    when "011" => spi1prescaler_var := 7;
                    when "100" => spi1prescaler_var := 15;
                    when "101" => spi1prescaler_var := 31;
                    when "110" => spi1prescaler_var := 63;
                    when "111" => spi1prescaler_var := 127;
                    when others => spi1prescaler_var  := 127;
                end case;

                -- If data register is read...
                -- Reading data register clears flags!
                if read_access_granted_second_cycle = '1' then
                    if reg_int = spi1data_addr then
                        -- Clear the received status bit
                        spi1.stat(3) <= '0';
                    end if;
                end if;
                
                -- Transmit/receive
                case spi1.state is
                    when idle =>
                        -- Clear receive buffer
                        spi1.rxbuffer <= (others => '0');
                        -- If start is active (data written)
                        if spi1.start = '1' then
                            -- Activate the NSS (slave select)
                            O_spi1nss <= '0';
                            spi1.state <= cssetup;
                            spi1.sck <= spi1.ctrl(2);
                            if spi1.ctrl(1) = '0' then
                                spi1.mosi <= spi1.txbuffer(31);
                            else
                                spi1.mosi <= spi1mosidefault;
                            end if;
                        else
                            spi1.mosi <= spi1mosidefault;
                        end if;
                        -- Load CS setup time before first clock
                        spi1.bittimer <= to_integer(unsigned(spi1.ctrl(27 downto 20)));
                    when cssetup =>
                        -- Wait CS setup time (+1 system clocks)
                        if spi1.bittimer > 0 then
                            spi1.bittimer <= spi1.bittimer - 1;
                        else
                            spi1.bittimer <= spi1prescaler_var;
                            spi1.state <= first;
                        end if;
                    when first =>
                        if spi1.bittimer > 0 then
                            spi1.bittimer <= spi1.bittimer - 1;
                        else
                            spi1.bittimer <= spi1prescaler_var;
                            spi1.state <= second;
                            spi1.sck <= not spi1.ctrl(2);
                            -- If CPHA is 0 ...
                            if spi1.ctrl(1) = '0' then
                                -- Clock in data from slave
                                spi1.rxbuffer <= spi1.rxbuffer(30 downto 0) & I_spi1miso;
                            else
                                -- CPHA = 1, write out data
                                spi1.txbuffer <= spi1.txbuffer(30 downto 0) & '0';
                                spi1.mosi <= spi1.txbuffer(31);
                            end if;
                        end if;
                    when second =>
                        if spi1.bittimer > 0 then
                            spi1.bittimer <= spi1.bittimer - 1;
                        else
                            spi1.bittimer <= spi1prescaler_var;
                            spi1.sck <= spi1.ctrl(2);
                            -- If CPHA is 0 ...
                            if spi1.ctrl(1) = '0' then
                                -- Clock out data
                                spi1.txbuffer <= spi1.txbuffer(30 downto 0) & '0';
                                spi1.mosi <= spi1.txbuffer(30);
                            else
                                -- Read in data from slave
                                spi1.rxbuffer <= spi1.rxbuffer(30 downto 0) & I_spi1miso;
                            end if;
                            -- Are still bits left to transmit?
                            if spi1.shiftcounter > 0 then
                                spi1.shiftcounter <= spi1.shiftcounter - 1;
                                spi1.state <= first;
                            else
                                -- All bits transferred
                                if spi1.ctrl(1) = '1' then
                                    -- CPHA = 1, half SPI clock leadout
                                    spi1.state <= leadout;
                                else
                                    -- Copy to data register
                                    spi1.data <= spi1.rxbuffer;
                                    -- Load CS hold time after last clock
                                    spi1.bittimer <= to_integer(unsigned(spi1.ctrl(19 downto 12)));
                                    -- Goto cshold
                                    spi1.state <= cshold;
                                end if;
                            end if;
                        end if;
                    when leadout =>
                        if spi1.bittimer > 0 then
                            spi1.bittimer <= spi1.bittimer - 1;
                        else
                            -- Load CS hold time after last clock
                            spi1.bittimer <= to_integer(unsigned(spi1.ctrl(19 downto 12)));
                            spi1.state <= cshold;
                        end if;
                        -- Copy to data register
                        spi1.data <= spi1.rxbuffer;
                    when cshold =>
                        -- Wait CS hold time
                        spi1.sck <= spi1.ctrl(2);
                        if spi1.bittimer > 0 then
                            spi1.bittimer <= spi1.bittimer - 1;
                        else
                            -- Disable NSS
                            O_spi1nss <= '1';
                            spi1.mosi <= spi1mosidefault;
                            -- Set the received status bit
                            spi1.stat(3) <= '1';
                            spi1.state <= idle;
                        end if;
                    when others => null;
                end case;
            end if; -- rising_edge
        end process;
        O_spi1sck <= spi1.sck;
        O_spi1mosi <= spi1.mosi;
    end generate;
    spi1gen_not : if not HAVE_SPI1 generate
        spi1.ctrl <= (others => '0');
        spi1.stat <= (others => '0');
        spi1.data <= (others =>'0');
        O_spi1sck <= 'Z';
        O_spi1mosi <= 'Z';
        O_spi1nss <= 'Z';
    end generate;


    --
    -- SPI2
    --
    spi2gen : if HAVE_SPI2 generate
        process (I_clk, I_areset) is
        --variable spi2txshiftcounter_var : integer range 0 to 31;
        variable spi2prescaler_v : integer range 0 to 255;
        begin
            -- Common resets et al.
            if I_areset = '1' then
                spi2.data <= (others => '0');
                spi2.ctrl <= (others => '0');
                spi2.stat <= (others => '0');
                spi2.start <= '0';
                spi2.state <= idle;
                spi2.txbuffer <= (others => '0');
                spi2.bittimer <= 0;
                spi2.shiftcounter <= 0;
                spi2.mosi <= spi2mosidefault;
                spi2.rxbuffer <= (others => '0');
                --spi2miso_sync <= '0';
                spi2.sck <= '0';
            elsif rising_edge(I_clk) then
                -- Default for start transmission
                spi2.start <= '0';
                -- Common register writes
                if write_access_granted = '1' then
                    if reg_int = spi2ctrl_addr then
                        -- A write to the control register
                        spi2.ctrl <= I_datain;
                        -- Set clock polarity
                        spi2.sck <= I_datain(2);
                    elsif reg_int = spi2stat_addr then
                        -- A write to the status register
                        spi2.stat <= I_datain;
                    elsif reg_int = spi2data_addr then
                        -- A write to the data register triggers a transmission
                        -- Signal start
                        spi2.start <= '1';
                        -- Load transmit buffer with 8/16/24/32 data bits
                        spi2.txbuffer <= (others => '0');
                        spi2.data <= (others => '0');
                        -- Load the desired bits to transfer
                        case spi2.ctrl(5 downto 4) is
                            when "00" =>   spi2.txbuffer(31 downto 24) <= I_datain(7 downto 0);
                                           spi2.shiftcounter <= 7;
                            when "01" =>   spi2.txbuffer(31 downto 16) <= I_datain(15 downto 0);
                                           spi2.shiftcounter <= 15;
                            when "10" =>   spi2.txbuffer(31 downto 8) <= I_datain(23 downto 0);
                                           spi2.shiftcounter <= 23;
                            when "11" =>   spi2.txbuffer <= I_datain;
                                           spi2.shiftcounter <= 31;
                            when others => spi2.txbuffer <= (others => '-');
                                           spi2.shiftcounter <= 0;
                        end case;
                        -- Signal that we are sending
                        spi2.stat(3) <= '0'; 
                    end if;
                end if;
                -- Zero out bits not needed
                spi2.ctrl(31 downto 11) <= (others => '0');
                spi2.ctrl(7 downto 6) <= (others => '0');
                spi2.ctrl(3) <= '0';
                spi2.ctrl(0) <= '0';
                spi2.stat(31 downto 4) <= (others => '0');
                spi2.stat(2 downto 0) <= (others =>'0');

                -- Calculate prescaler, 2 to 256 in powers of 2
                case spi2.ctrl(10 downto 8) is
                    when "000" =>  spi2prescaler_v := 0;
                    when "001" =>  spi2prescaler_v := 1;
                    when "010" =>  spi2prescaler_v := 3;
                    when "011" =>  spi2prescaler_v := 7;
                    when "100" =>  spi2prescaler_v := 15;
                    when "101" =>  spi2prescaler_v := 31;
                    when "110" =>  spi2prescaler_v := 63;
                    when "111" =>  spi2prescaler_v := 127;
                    when others => spi2prescaler_v  := 127;
                end case;

                -- If data register is read...
                -- Reading data register clears flags!
                if read_access_granted_second_cycle = '1' then
                    if reg_int = spi2data_addr then
                        -- Clear the received status bit
                        spi2.stat(3) <= '0';
                    end if;
                end if;
                
                -- Transmit/receive
                case spi2.state is
                    when idle =>
                        -- Clear receive buffer
                        spi2.rxbuffer <= (others => '0');
                        -- Load prescaler value
                        spi2.bittimer <= spi2prescaler_v;
                        -- If start is active (data written)
                        if spi2.start = '1' then
                            spi2.state <= first;
                            spi2.sck <= spi2.ctrl(2);
                            if spi2.ctrl(1) = '0' then
                                spi2.mosi <= spi2.txbuffer(31);
                            else
                                -- CPHA = 1, write out data
                                spi2.txbuffer <= spi2.txbuffer(30 downto 0) & '0';
                                spi2.mosi <= spi2.txbuffer(31);
                                spi2.sck <= not spi2.ctrl(2);
                                spi2.state <= second;
                            end if;
                        else
                            spi2.mosi <= spi2mosidefault;
                        end if;
                    when first =>
                        if spi2.bittimer > 0 then
                            spi2.bittimer <= spi2.bittimer - 1;
                        else
                            spi2.bittimer <= spi2prescaler_v;
                            spi2.state <= second;
                            spi2.sck <= not spi2.ctrl(2);
                            if spi2.ctrl(1) = '0' then
                                -- CPHA = 0, clock in data from slave
                                spi2.rxbuffer <= spi2.rxbuffer(30 downto 0) & I_spi2miso;
                            else
                                -- CPHA = 1, write out data
                                spi2.txbuffer <= spi2.txbuffer(30 downto 0) & '0';
                                spi2.mosi <= spi2.txbuffer(31);
                            end if;
                        end if;
                    when second =>
                        if spi2.bittimer > 0 then
                            spi2.bittimer <= spi2.bittimer - 1;
                        else
                            spi2.bittimer <= spi2prescaler_v;
                            spi2.sck <= spi2.ctrl(2);
                            if spi2.ctrl(1) = '0' then
                                -- If CPHA is 0, clock out data
                                spi2.txbuffer <= spi2.txbuffer(30 downto 0) & '0';
                                -- Must be spi2buffer(30) because data is not yet shifted
                                spi2.mosi <= spi2.txbuffer(30);
                            else
                                -- If CPHA = 1, read in data from slave
                                spi2.rxbuffer <= spi2.rxbuffer(30 downto 0) & I_spi2miso;
                            end if;
                            -- Are still bits left to transmit?
                            if spi2.shiftcounter > 0 then
                                spi2.shiftcounter <= spi2.shiftcounter - 1;
                                spi2.state <= first;
                            else
                                -- All bits transferred
                                if spi2.ctrl(1) = '1' then
                                    -- CPHA = 1, half SPI clock leadout
                                    spi2.state <= leadout;
                                else
                                    -- CPHA = 0, no leadout, goto idle
                                    spi2.sck <= spi2.ctrl(2);
                                    spi2.stat(3) <= '1';
                                    spi2.mosi <= spi2mosidefault;
                                    spi2.state <= idle;
                                    -- Copy to data register
                                    spi2.data <= spi2.rxbuffer;
                                end if;
                            end if;
                        end if;
                    when leadout =>
                        -- Hold the data half SPI clock cycle
                        if spi2.bittimer > 0 then
                            spi2.bittimer <= spi2.bittimer - 1;
                        else
                            spi2.sck <= spi2.ctrl(2);
                            spi2.stat(3) <= '1';
                            spi2.mosi <= spi2mosidefault;
                            spi2.state <= idle;
                        end if;
                        -- Copy to data register
                        spi2.data <= spi2.rxbuffer;
                when others => null;
                end case;
            end if; -- rising_edge
        end process;
        O_spi2sck <= spi2.sck;
        O_spi2mosi <= spi2.mosi;
    end generate;
    spi2gen_not : if not HAVE_SPI2 generate
        spi2.ctrl <= (others => '0');
        spi2.stat <= (others => '0');
        spi2.data <= (others =>'0');
        O_spi2sck <= 'Z';
        O_spi2mosi <= 'Z';
    end generate;

    
    --
    -- TIMER1 - a very simple timer
    --
    timer1gen : if HAVE_TIMER1 generate
        process (I_clk, I_areset) is
        begin
            if I_areset = '1' then
                timer1.ctrl <= (others => '0');
                timer1.stat <= (others => '0');
                timer1.cntr <= (others => '0');
                timer1.cmpt <= (others => '0');
            elsif rising_edge(I_clk) then
                if write_access_granted = '1' then
                    -- Write Timer Control Register
                    if reg_int = timer1ctrl_addr then
                        timer1.ctrl <= I_datain;
                    end if;
                    -- Write Timer Status Register
                    if reg_int = timer1stat_addr then
                        timer1.stat <= I_datain;
                    end if;
                    -- Write Timer Counter Register
                    if reg_int = timer1cntr_addr then
                        timer1.cntr <= I_datain;
                    end if;
                    -- Write Timer Compare Register
                    if reg_int = timer1cmpt_addr then
                        timer1.cmpt <= I_datain;
                    end if;
                end if;
                -- Set unused bits to 0
                timer1.ctrl(31 downto 12) <= (others => '0');
                timer1.stat(31 downto 12) <= (others => '0');
                
                -- If timer is enabled....
                if timer1.ctrl(0) = '1' then
                    -- If we hit the Compare Register T...
                    if timer1.cntr >= timer1.cmpt then
                        -- Reload Counter Register
                        timer1.cntr <= (others => '0');
                        -- Signal hit
                        timer1.stat(4) <= '1';
                    else
                        -- else, increment the Counter Register
                        timer1.cntr <= std_logic_vector(unsigned(timer1.cntr) + 1);
                    end if;
                end if;
            end if;
        end process;
    end generate;
    timer1gen_not : if not HAVE_TIMER1 generate
        timer1.ctrl <= (others => '0');
        timer1.stat <= (others => '0');
        timer1.cntr <= (others => '0');
        timer1.cmpt <= (others => '0');
    end generate;

    --
    -- TIMER2 - a more elaborate timer
    --
    timer2gen : if HAVE_TIMER2 generate
        process (I_clk, I_areset) is
        begin
            if I_areset = '1' then
                -- The I/O registers
                timer2.ctrl <= (others => '0');
                timer2.stat <= (others => '0');
                timer2.cntr <= (others => '0');
                timer2.cmpt <= (others => '0');
                timer2.prsc <= (others => '0');
                timer2.cmpa <= (others => '0');
                timer2.cmpb <= (others => '0');
                timer2.cmpc <= (others => '0');
                -- The internal prescaler
                timer2.prescaler <= (others => '0');
                -- The shadow registers
                timer2.prscshadow <= (others => '0');
                timer2.cmptshadow <= (others => '0');
                timer2.cmpashadow <= (others => '0');
                timer2.cmpbshadow <= (others => '0');
                timer2.cmpcshadow <= (others => '0');
                -- The OC outputs
                timer2.oct <= '0';
                timer2.oca <= '0';
                timer2.ocb <= '0';
                timer2.occ <= '0';
                -- The IC synchronizers
                timer2.icasync <= (others => '0');
                timer2.icbsync <= (others => '0');
                timer2.iccsync <= (others => '0');
            elsif rising_edge(I_clk) then
                if write_access_granted = '1' then
                    -- Write Timer Control Register
                    if reg_int = timer2ctrl_addr then
                        -- Check if one or more FOC bits are set
                        -- If so, the data is NOT copied to the CTRL register
                        -- and the MODE bits indicate the FOC action
                        if I_datain(31 downto 28) /= "0000" then
                            -- FOCT
                            if I_datain(28) = '1' then
                                case I_datain(14 downto 12) is
                                    when "001" => timer2.oct <= not timer2.oct;
                                    when "010" => timer2.oct <= '1';
                                    when "011" => timer2.oct <= '0';
                                    when others => null;
                                end case;
                            end if;
                            -- FOCA
                            if I_datain(29) = '1' then
                                case I_datain(18 downto 16) is
                                    when "001" => timer2.oca <= not timer2.oca;
                                    when "010" => timer2.oca <= '1';
                                    when "011" => timer2.oca <= '0';
                                    when others => null;
                                end case;
                            end if;
                            -- FOCB
                            if I_datain(30) = '1' then
                                case I_datain(22 downto 20) is
                                    when "001" => timer2.ocb <= not timer2.ocb;
                                    when "010" => timer2.ocb <= '1';
                                    when "011" => timer2.ocb <= '0';
                                    when others => null;
                                end case;
                            end if;
                            -- FOCC
                            if I_datain(31) = '1' then
                                case I_datain(26 downto 24) is
                                    when "001" => timer2.occ <= not timer2.occ;
                                    when "010" => timer2.occ <= '1';
                                    when "011" => timer2.occ <= '0';
                                    when others => null;
                                end case;
                            end if;
                        else
                            -- No FOC bits set, so ...
                            -- Copy to CTRL register
                            timer2.ctrl <= I_datain;
                            -- Set the signal phase
                            timer2.oct <= I_datain(15);
                            timer2.oca <= I_datain(19);
                            timer2.ocb <= I_datain(23);
                            timer2.occ <= I_datain(27);
                            -- If the CMPA register is all zero and we start, then
                            -- set the output compare immediate, but don't flag it
                            if timer2.cmpa = x"00000000" and I_datain(0) = '1' then
                                if I_datain(18 downto 16) = "001" then
                                    timer2.oca <= not I_datain(19);
                                elsif I_datain(18 downto 16) = "010" and I_datain(0) = '1' then
                                    timer2.oca <= not I_datain(19);
                                elsif I_datain(18 downto 16) = "011" and I_datain(0) = '1' then
                                    timer2.oca <= I_datain(19);
                                end if;
                            end if;
                            -- If the CMPB register is all zero and we start, then
                            -- set the output compare immediate, but don't flag it
                            if timer2.cmpb = x"00000000" and I_datain(0) = '1' then
                                if I_datain(22 downto 20) = "001" then
                                    timer2.ocb <= not I_datain(23);
                                elsif I_datain(22 downto 20) = "010" and I_datain(0) = '1' then
                                    timer2.ocb <= not I_datain(23);
                                elsif I_datain(22 downto 20) = "011" and I_datain(0) = '1' then
                                    timer2.ocb <= I_datain(23);
                                end if;
                            end if;
                            -- If the CMPC register is all zero and we start, then
                            -- set the output compare immediate, but don't flag it
                            if timer2.cmpc = x"00000000" and I_datain(0) = '1' then
                                if I_datain(26 downto 24) = "001" then
                                    timer2.occ <= not I_datain(27);
                                elsif I_datain(26 downto 24) = "010" and I_datain(0) = '1' then
                                    timer2.occ <= not I_datain(27);
                                elsif I_datain(26 downto 24) = "011" and I_datain(0) = '1' then
                                    timer2.occ <= I_datain(27);
                                end if;
                            end if;
                        end if;
                    end if;
                    -- Write Timer Status Register
                    if reg_int = timer2stat_addr then
                        timer2.stat <= I_datain;
                    end if;
                    -- Write Timer Counter Register
                    if reg_int = timer2cntr_addr then
                        timer2.cntr <= I_datain;
                    end if;
                    -- Write Timer Compare T Register
                    if reg_int = timer2cmpt_addr then
                        timer2.cmpt <= I_datain;
                        -- If the timer is stopped or preload is off, directly write the shadow register
                        if timer2.ctrl(0) = '0' or timer2.ctrl(8) = '0' then
                            timer2.cmptshadow <= I_datain;
                        end if;
                    end if;
                    -- Write Prescaler Register
                    if reg_int = timer2prsc_addr then
                        timer2.prsc <= I_datain;
                        -- If the timer is stopped, directly write the shadow register
                        if timer2.ctrl(0) = '0' then
                            timer2.prscshadow <= I_datain;
                        end if;
                        -- Reset internal prescaler
                        timer2.prescaler <= (others => '0');
                    end if;
                    -- Write Timer Compare A Register
                    if reg_int = timer2cmpa_addr then
                        timer2.cmpa <= I_datain;
                        -- If the timer is stopped or preload is off, directly write the shadow register
                        if timer2.ctrl(0) = '0' or timer2.ctrl(9) = '0' then
                            timer2.cmpashadow <= I_datain;
                        end if;
                    end if;
                    -- Write Timer Compare B Register
                    if reg_int = timer2cmpb_addr then
                        timer2.cmpb <= I_datain;
                        -- If the timer is stopped or preload is off, directly write the shadow register
                        if timer2.ctrl(0) = '0' or timer2.ctrl(10) = '0' then
                            timer2.cmpbshadow <= I_datain;
                        end if;
                    end if;
                    -- Write Timer Compare C Register
                    if reg_int = timer2cmpc_addr then
                        timer2.cmpc <= I_datain;
                        -- If the timer is stopped or preload is off, directly write the shadow register
                        if timer2.ctrl(0) = '0' or timer2.ctrl(11) = '0' then
                            timer2.cmpcshadow <= I_datain;
                        end if;
                    end if;
                end if;
                -- Set unused bits to 0 for CTRL and STAT
                timer2.ctrl(31 downto 28) <= (others => '0');
                timer2.stat(31 downto 12) <= (others => '0');
                
                -- If timer is enabled....
                if timer2.ctrl(0) = '1' then
                    -- If internal prescaler at end...
                    if timer2.prescaler >= timer2.prscshadow then
                        -- Wrap internal prescaler
                        timer2.prescaler <= (others => '0');
                        -- If we hit the Compare Register T...
                        if timer2.cntr >= timer2.cmptshadow then
                            -- Clear Counter Register
                            timer2.cntr <= (others => '0');
                            -- Signal hit
                            timer2.stat(4) <= '1';
                            -- Toggle OCT, or not
                            case timer2.ctrl(14 downto 12) is
                                when "000" => timer2.oct <= '0'; -- off
                                when "001" => timer2.oct <= not timer2.oct; -- toggle
                                when "010" => timer2.oct <= not timer2.ctrl(15); -- invert PHAT
                                when "011" => timer2.oct <= timer2.ctrl(15); -- write PHAT
                                -- Others not allowed, as T does not have PWM mode
                                when others => timer2.oct <= '0';
                            end case;
                            -- If we have a one-shot, disable timer
                            if timer2.ctrl(3) = '1' then
                                timer2.ctrl(0) <= '0';
                                timer2.prescaler <= (others => '0');
                                --timer2cntr_int <= (others => '0');
                            end if;
                        else
                            -- If we are at the last step - 1 ...
                            if timer2.cntr = std_logic_vector(unsigned(timer2.cmptshadow)-1) then
                                -- Load PRSC shadow register
                                timer2.prscshadow <= timer2.prsc;
                                -- Load CMPT shadow register
                                timer2.cmptshadow <= timer2.cmpt;
                                -- Load CMPA shadow register
                                timer2.cmpashadow <= timer2.cmpa;
                                -- Load CMPB shadow register
                                timer2.cmpbshadow <= timer2.cmpb;
                                -- Load CMPC shadow register
                                timer2.cmpcshadow <= timer2.cmpc;
                            end if;
                            -- else, increment the Counter Register
                            timer2.cntr <= std_logic_vector(unsigned(timer2.cntr) + 1);
                        end if;
                    else
                        timer2.prescaler <= std_logic_vector(unsigned(timer2.prescaler) + 1);
                    end if;
                    -- If we are at the end of prescale counting
                    if timer2.prescaler >= timer2.prscshadow then
                        -- Sync the IC inputs
                        timer2.icasync <= timer2.icasync(1 downto 0) & IO_timer2icoca;
                        timer2.icbsync <= timer2.icbsync(1 downto 0) & IO_timer2icocb;
                        timer2.iccsync <= timer2.iccsync(1 downto 0) & IO_timer2icocc;
                    
                        -- Check CMPA for mode
                        case timer2.ctrl(18 downto 16) is
                            -- 000 = do nothing
                            when "000" => timer2.oca <= '0';
                            -- 001 = toggle on compare match
                            when "001" =>
                                if timer2.cmpashadow = x"00000000" and timer2.cntr = timer2.cmptshadow then
                                    timer2.oca <= not timer2.oca;
                                    timer2.stat(5) <= '1';
                                elsif timer2.cntr = std_logic_vector(unsigned(timer2.cmpashadow)-1) then
                                    timer2.oca <= not timer2.oca;
                                    timer2.stat(5) <= '1';
                                end if;
                            -- 010 = activate on compare match, invert PHAA
                            when "010" =>
                                if timer2.cmpashadow = x"00000000" and timer2.cntr = timer2.cmptshadow then
                                    timer2.oca <= not timer2.ctrl(19);
                                    timer2.stat(5) <= '1';
                                elsif timer2.cntr = std_logic_vector(unsigned(timer2.cmpashadow)-1) then
                                    timer2.oca <= not timer2.ctrl(19);
                                    timer2.stat(5) <= '1';
                                end if;
                            -- 011 = deactivate on compare match, write PHAA
                            when "011" =>
                                if timer2.cmpashadow = x"00000000" and timer2.cntr = timer2.cmptshadow then
                                    timer2.oca <= timer2.ctrl(19);
                                    timer2.stat(5) <= '1';
                                elsif timer2.cntr = std_logic_vector(unsigned(timer2.cmpashadow)-1) then
                                    timer2.oca <= timer2.ctrl(19);
                                    timer2.stat(5) <= '1';
                                end if;
                            -- 100 = edge aligned PWM
                            when "100" =>
                                if timer2.cmpashadow = x"00000000" then
                                    timer2.oca <= timer2.ctrl(19);
                                elsif timer2.cntr < std_logic_vector(unsigned(timer2.cmpashadow)-1) or (timer2.cntr = timer2.cmptshadow and timer2.ctrl(3) = '0') then
                                    timer2.oca <= not timer2.ctrl(19);
                                else
                                    timer2.oca <= timer2.ctrl(19);
                                end if;
                                if timer2.cntr = std_logic_vector(unsigned(timer2.cmpashadow)-1) then
                                    timer2.stat(5) <= '1';
                                end if;
                            -- 110 - positive edge detected
                            when "110" =>
                                if timer2.icasync(2 downto 1) = "01" then
                                    -- Copy CNTR to CMPA register and raise interrupt
                                    timer2.cmpa <= timer2.cntr;
                                    timer2.stat(5) <= '1';
                                end if;
                            -- 111 - negative edge detected
                            when "111" =>
                                if timer2.icasync(2 downto 1) = "10" then
                                    -- Copy CNTR to CMPA register and raise interrupt
                                    timer2.cmpa <= timer2.cntr;
                                    timer2.stat(5) <= '1';
                                end if;
                            -- Others not allowed
                            when others => timer2.oca <= '0';
                        end case;
                        -- Check CMPB for mode
                    case timer2.ctrl(22 downto 20) is
                        -- 000 = do nothing
                        when "000" => timer2.ocb <= '0';
                        -- 001 = toggle on compare match
                        when "001" =>
                            if timer2.cmpbshadow = x"00000000" and timer2.cntr = timer2.cmptshadow then
                                timer2.ocb <= not timer2.ocb;
                                timer2.stat(6) <= '1';
                            elsif timer2.cntr = std_logic_vector(unsigned(timer2.cmpbshadow)-1) then
                                timer2.ocb <= not timer2.ocb;
                                timer2.stat(6) <= '1';
                            end if;
                        -- 010 = activate on compare match, invert PHAB
                        when "010" =>
                            if timer2.cmpbshadow = x"00000000" and timer2.cntr = timer2.cmptshadow then
                                timer2.ocb <= not timer2.ctrl(23);
                                timer2.stat(6) <= '1';
                            elsif timer2.cntr = std_logic_vector(unsigned(timer2.cmpbshadow)-1) then
                                timer2.ocb <= not timer2.ctrl(23);
                                timer2.stat(6) <= '1';
                            end if;
                        -- 011 = deactivate on compare match, write PHAB
                        when "011" =>
                            if timer2.cmpbshadow = x"00000000" and timer2.cntr = timer2.cmptshadow then
                                timer2.ocb <= timer2.ctrl(23);
                                timer2.stat(6) <= '1';
                            elsif timer2.cntr = std_logic_vector(unsigned(timer2.cmpbshadow)-1) then
                                timer2.ocb <= timer2.ctrl(23);
                                timer2.stat(6) <= '1';
                            end if;
                        -- 100 = edge aligned PWM
                        when "100" =>
                            if timer2.cmpbshadow = x"00000000" then
                                timer2.ocb <= timer2.ctrl(23);
                            elsif timer2.cntr < std_logic_vector(unsigned(timer2.cmpbshadow)-1) or (timer2.cntr = timer2.cmptshadow and timer2.ctrl(3) = '0') then
                                timer2.ocb <= not timer2.ctrl(23);
                            else
                                timer2.ocb <= timer2.ctrl(23);
                            end if;
                            if timer2.cntr = std_logic_vector(unsigned(timer2.cmpbshadow)-1) then
                                timer2.stat(6) <= '1';
                            end if;
                        -- 110 - positive edge detected
                        when "110" =>
                            if timer2.icbsync(2 downto 1) = "01" then
                                -- Copy CNTR to CMPB register and raise interrupt
                                timer2.cmpb <= timer2.cntr;
                                timer2.stat(6) <= '1';
                            end if;
                        -- 111 - negative edge detected
                        when "111" =>
                            if timer2.icbsync(2 downto 1) = "10" then
                                -- Copy CNTR to CMPB register and raise interrupt
                                timer2.cmpb <= timer2.cntr;
                                timer2.stat(6) <= '1';
                            end if;
                        when others => timer2.ocb <= '0';
                    end case;
                        -- Check CMPC for mode
                        case timer2.ctrl(26 downto 24) is
                            -- 000 = do nothing
                            when "000" => timer2.occ <= '0';
                            -- 001 = toggle on compare match
                            when "001" =>
                                if timer2.cmpcshadow = x"00000000" and timer2.cntr = timer2.cmptshadow then
                                    timer2.occ <= not timer2.occ;
                                    timer2.stat(7) <= '1';
                                elsif timer2.cntr = std_logic_vector(unsigned(timer2.cmpcshadow)-1) then
                                    timer2.occ <= not timer2.occ;
                                    timer2.stat(7) <= '1';
                                end if;
                            -- 010 = activate on compare match, invert PHAC
                            when "010" =>
                                if timer2.cmpcshadow = x"00000000" and timer2.cntr = timer2.cmptshadow then
                                    timer2.occ <= not timer2.ctrl(27);
                                    timer2.stat(7) <= '1';
                                elsif timer2.cntr = std_logic_vector(unsigned(timer2.cmpcshadow)-1) then
                                    timer2.occ <= not timer2.ctrl(27);
                                    timer2.stat(7) <= '1';
                                end if;
                            -- 011 = deactivate on compare match, write PHAC
                            when "011" =>
                                if timer2.cmpcshadow = x"00000000" and timer2.cntr = timer2.cmptshadow then
                                    timer2.occ <= timer2.ctrl(27);
                                    timer2.stat(7) <= '1';
                                elsif timer2.cntr = std_logic_vector(unsigned(timer2.cmpcshadow)-1) then
                                    timer2.occ <= timer2.ctrl(27);
                                    timer2.stat(7) <= '1';
                                end if;
                            -- 100 = edge aligned PWM
                            when "100" =>
                                if timer2.cmpcshadow = x"00000000" then
                                    timer2.occ <= timer2.ctrl(27);
                                elsif timer2.cntr < std_logic_vector(unsigned(timer2.cmpcshadow)-1) or (timer2.cntr = timer2.cmptshadow and timer2.ctrl(3) = '0') then
                                    timer2.occ <= not timer2.ctrl(27);
                                else
                                    timer2.occ <= timer2.ctrl(27);
                                end if;
                                if timer2.cntr = std_logic_vector(unsigned(timer2.cmpcshadow)-1) then
                                    timer2.stat(7) <= '1';
                                end if;
                            -- 110 - positive edge detected
                            when "110" =>
                                if timer2.iccsync(2 downto 1) = "01" then
                                    -- Copy CNTR to CMPC register and raise interrupt
                                    timer2.cmpc <= timer2.cntr;
                                    timer2.stat(7) <= '1';
                                end if;
                            -- 111 - negative edge detected
                            when "111" =>
                                if timer2.iccsync(2 downto 1) = "10" then
                                    -- Copy CNTR to CMPC register and raise interrupt
                                    timer2.cmpc <= timer2.cntr;
                                    timer2.stat(7) <= '1';
                                end if;
                            when others => timer2.occ <= '0';
                        end case;
                    end if;
                else
                end if;
                -- Set unused bits, all counter registers are 16 bits.
                timer2.cntr(31 downto 16) <= (others => '0');
                timer2.cmpt(31 downto 16) <= (others => '0');
                timer2.prsc(31 downto 16) <= (others => '0');
                timer2.cmpa(31 downto 16) <= (others => '0');
                timer2.cmpb(31 downto 16) <= (others => '0');
                timer2.cmpc(31 downto 16) <= (others => '0');
                timer2.prescaler(31 downto 16) <= (others => '0');
                timer2.prscshadow(31 downto 16) <= (others => '0');
                timer2.cmptshadow(31 downto 16) <= (others => '0');
                timer2.cmpashadow(31 downto 16) <= (others => '0');
                timer2.cmpbshadow(31 downto 16) <= (others => '0');
                timer2.cmpcshadow(31 downto 16) <= (others => '0');
            end if;
        end process;
        -- Generate Output Enabled
        timer2.ocaen <= '1' when timer2.ctrl(18 downto 16) = "001" or
                                    timer2.ctrl(18 downto 16) = "010" or
                                    timer2.ctrl(18 downto 16) = "011" or
                                    timer2.ctrl(18 downto 16) = "100"
                               else '0';
        timer2.ocben <= '1' when timer2.ctrl(22 downto 20) = "001" or
                                    timer2.ctrl(22 downto 20) = "010" or
                                    timer2.ctrl(22 downto 20) = "011" or
                                    timer2.ctrl(22 downto 20) = "100"
                               else '0';
        timer2.occen <= '1' when timer2.ctrl(26 downto 24) = "001" or
                                    timer2.ctrl(26 downto 24) = "010" or
                                    timer2.ctrl(26 downto 24) = "011" or
                                    timer2.ctrl(26 downto 24) = "100"
                               else '0';
        -- Output the Output Compare match
        O_timer2oct <= timer2.oct;
        IO_timer2icoca <= timer2.oca when timer2.ocaen = '1' else 'Z';
        IO_timer2icocb <= timer2.ocb when timer2.ocben = '1' else 'Z';
        IO_timer2icocc <= timer2.occ when timer2.occen = '1' else 'Z';
    end generate;
    timer2gen_not : if not HAVE_TIMER2 generate
        timer2.ctrl <= (others => '0');
        timer2.stat <= (others => '0');
        timer2.cntr <= (others => '0');
        timer2.cmpt <= (others => '0');
        timer2.prsc <= (others => '0');
        timer2.cmpa <= (others => '0');
        timer2.cmpb <= (others => '0');
        timer2.cmpc <= (others => '0');
        O_timer2oct <= 'Z';
        IO_timer2icoca <= 'Z';
        IO_timer2icocb <= 'Z';
        IO_timer2icocc <= 'Z';
    end generate;

    
    --
    -- RISC-V Machine Software Interrupt (MSI)
    --
    process (I_clk, I_areset) is
    begin
        if I_areset = '1' then
            msi.trig(0) <= '0';
        elsif rising_edge(I_clk) then
            if write_access_granted = '1' then
                -- Set trigger bit
                if reg_int = msitrig_addr then
                    msi.trig(0) <= I_datain(0);
                end if;
            end if;
        end if;
    end process;
    msi.trig(31 downto 1) <= (others => '0');
    
    
    --
    -- RISC-V system timer TIME and TIMECMP
    -- These registers are memory mapped
    --
    process (I_clk, I_areset, mtime) is
    variable mtime_v : unsigned(63 downto 0);
    variable mtimecmp_v : unsigned(63 downto 0);
    variable prescaler_v : integer range 0 to SYSTEM_FREQUENCY/CLOCK_FREQUENCY-1;
    begin
        if I_areset = '1' then
            mtime_v := (others => '0');
            mtimecmp_v := (others => '0');
            prescaler_v := 0;
        elsif rising_edge(I_clk) then
            if write_access_granted = '1' then
                -- Load time (low 32 bits)
                if reg_int = mtime_addr then
                    mtime_v(31 downto 0) := unsigned(I_datain);
                end if;
                -- Load timeh (high 32 bits)
                if reg_int = mtimeh_addr then
                    mtime_v(63 downto 32) := unsigned(I_datain);
                end if;
                -- Load compare register (low 32 bits)
                if reg_int = mtimecmp_addr then
                    mtimecmp_v(31 downto 0) := unsigned(I_datain);
                end if;
                -- Load compare register (high 32 bits)
                if reg_int = mtimecmph_addr then
                    mtimecmp_v(63 downto 32) := unsigned(I_datain);
                end if;
            end if;
            -- Update system timer
            if prescaler_v = SYSTEM_FREQUENCY/CLOCK_FREQUENCY-1 then
                prescaler_v := 0;
                mtime_v := mtime_v + 1;
            else
                prescaler_v := prescaler_v + 1;
            end if;
        end if;
        mtime.mtime <= std_logic_vector(mtime_v(31 downto 0));
        mtime.mtimeh <= std_logic_vector(mtime_v(63 downto 32));
        mtime.mtimecmp <= std_logic_vector(mtimecmp_v(31 downto 0));
        mtime.mtimecmph <= std_logic_vector(mtimecmp_v(63 downto 32));
        -- If compare register >= time register, assert interrupt
        if mtime_v >= mtimecmp_v then
            O_intrio(INTR_PRIO_MTIME) <= '1';
        else
            O_intrio(INTR_PRIO_MTIME) <= '0';
        end if;
        O_mtime <= mtime.mtime;
        O_mtimeh <= mtime.mtimeh;
    end process;
    
    --
    -- Interrupt generation
    --

    process (spi1, i2c1, i2c2, timer2, timer1, uart1, gpioa, msi) is
    begin
       -- Default all interrupts to 0.
        O_intrio(31 downto 8) <= (others => '0');
       -- System Timer is handled by timer hardware
        O_intrio(6 downto 0) <= (others => '0');

        -- SPI1 transmit complete interrupt
        if spi1.ctrl(3) = '1' and spi1.stat(3) = '1' then
            O_intrio(INTR_PRIO_SPI1) <= '1';
        end if;
        -- I2C1 transmit interrupt.
        if i2c1.ctrl(3) = '1' and i2c1.stat(3) = '1' then
            O_intrio(INTR_PRIO_I2C1) <= '1';
        end if;
        -- I2C2 transmit interrupt.
        if i2c2.ctrl(3) = '1' and i2c2.stat(3) = '1' then
            O_intrio(INTR_PRIO_I2C2) <= '1';
        end if;
        -- TIMER2 compare match T/A/B/C interrupt
        if (timer2.ctrl(4) = '1' and timer2.stat(4) = '1') or
           (timer2.ctrl(5) = '1' and timer2.stat(5) = '1') or
           (timer2.ctrl(6) = '1' and timer2.stat(6) = '1') or
           (timer2.ctrl(7) = '1' and timer2.stat(7) = '1') then
            O_intrio(INTR_PRIO_TIMER2) <= '1';
        end if;
        -- UART1 receive or transmit interrupt. Software must determine if it was
        -- receive or transmit or both
        if (uart1.stat(4) = '1' and uart1.ctrl(7) = '1') or
           (uart1.stat(2) = '1' and uart1.ctrl(6) = '1') then
            O_intrio(INTR_PRIO_UART1) <= '1';
        end if;
        -- TIMER1 compare match interrupt
        if timer1.ctrl(4) = '1' and timer1.stat(4) = '1' then
            O_intrio(INTR_PRIO_TIMER1) <= '1';
        end if;
        -- EXTI external input interrupt
        if gpioa.exts(0) = '1' then
            O_intrio(INTR_PRIO_EXTI) <= '1';
        end if;
        --
        if msi.trig(0) = '1' then
            O_intrio(INTR_PRIO_MSI) <= '1';
        end if;
    end process;


    -- This process determines if a side effect of reading a register may proceed.
    -- Side effect: reading a data register (e.g. UART1, SPI1/2, I2C) clears flags
    -- in the status register, but only if the read (LOAD) is not interrupted by
    -- an assertion of an interrupt request.
    process (I_clk, I_areset) is
    begin
        if I_areset = '1' then
            read_access_granted_ff <= '0';
        elsif rising_edge(I_clk) then
            if read_access_granted = '1' and read_access_granted_ff = '0' then
                read_access_granted_ff <= '1';
            else
                read_access_granted_ff <= '0';
            end if;
        end if;
    end process;
    read_access_granted_second_cycle <= read_access_granted_ff and read_access_granted;

        
    -- Generate I/O ready signal for reads and writes
    -- This is faster than using read_access_granted and write_access_granted
    process (I_clk, I_areset, I_csio, I_wren) is
    begin
        if I_areset = '1' then
            readready <= '0';
        elsif rising_edge(I_clk) then
            if readready = '1' then
                readready <= '0';
            elsif I_csio = '1' and I_wren = '0' then
                readready <= '1';
            else
                readready <= '0';
            end if;
        end if;

    end process;

    -- Fuse read ready and write ready
    O_memready <= readready  or (I_csio and I_wren and boolean_to_std_logic(not HAVE_FAST_STORE));
   
    -- Only for view in the simulator 
-- synthesis translate_off
    io_alt <= (
         0 => gpioa.pin,
         1 => gpioa.pout,
         -- 2 - 5 not used
         6 => gpioa.extc,
         7 => gpioa.exts,
         8 => uart1.ctrl,
         9 => uart1.stat,
        10 => uart1.data,
        11 => uart1.baud,
        -- 12 - 15 not used
        16 => i2c1.ctrl,
        17 => i2c1.stat,
        18 => i2c1.data,
        -- 19 not used
        20 => i2c2.ctrl,
        21 => i2c2.stat,
        22 => i2c2.data,
        -- 23 not used
        24 => spi1.ctrl,
        25 => spi1.stat,
        26 => spi1.data,
        -- 27 not used
        28 => spi2.ctrl,
        29 => spi2.stat,
        30 => spi2.data,
        -- 31 not used
        32 => timer1.ctrl,
        33 => timer1.stat,
        34 => timer1.cntr,
        35 => timer1.cmpt,
        -- 36 - 39 not used
        40 => timer2.ctrl,
        41 => timer2.stat,
        42 => timer2.cntr,
        43 => timer2.cmpt,
        44 => timer2.prsc,
        45 => timer2.cmpa,
        46 => timer2.cmpb,
        47 => timer2.cmpc,
        -- 48 - 58 not used
        59 => msi.trig,
        60 => mtime.mtime,
        61 => mtime.mtimeh,
        62 => mtime.mtimecmp,
        63 => mtime.mtimecmph,
        others => (others => 'X')
       );
-- synthesis translate_on
    
end architecture rtl;
